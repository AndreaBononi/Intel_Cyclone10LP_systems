//__ACDS_USER_COMMENT__ (C) 2001-2023 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
//__ACDS_USER_COMMENT__ ACDS 22.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
GXarB8PdlOqLa+xm5vExLiiUfu6H9rZbqbJc+wEgC/cwD4qCchBh4QsdTq6y+HyU15llaqzD8uWv
d7OvGqdykQDyzColZlvpITS6DX0o4kq+XtPFJsbXa4I4ZC/g2PCc1JYWYC5G0gceLulA00Igyzrq
/sj4KQqZ1Wj5ZWB2J1SkkKbFLGIiDb8pqSsUX+37R37CvA1WuwpRKZB+eWokl3d7tD1PecEUlWdG
siEmDvGmbgfxYVDMoJrJHZXKaG/ioID4wAubObK15Phvtw0nirF90fKX0SsgDvATlfwMpnGh2WRC
hzn5Bu9pTHkaVAiHkBeK/Tzuo2/NVnoZAExRCg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12256)
XW5LXafsQKsB6JfZltSqR94cmmYNClrIVRHzYXSYnj2dZ/sszb7Es0gdyOMp8DlRXmOqBDART3M2
tMHvs90GFuiHJUtMJP1/iYl2o8BV1rvvMQKHS0Er7hoA7uVcffZW4YVa4tRXR/k6d0MPsfTn0VO4
zdHxXYcTjEGZkQX5M8rNFVq0UkCWeeoee4pos0imy/HBbu/xUpEnTgPZ+rkdIvRs42YjuD04dQKH
HBRWbMtFzm2OIuQknS7Kj8GtqPbK7UoCvM5/wpZP29Yp0sK57XnN2VJ1PDSYJbSk5V3G3jpUbChu
G6Imdf1GZ9OgeaYnLBl81Tl0Iq8Bnp4O1QNtPVTp+mKnEc6Jwo6hrndhgFbmF6yQpn9Cm9D/70HR
5/QQNn9WeoyHLZLtP7IF9oNiz8xR5EsxTDBYhEU5kNQBUUzzFf6yrD5biP2tkihoibBhh/XsHbTP
4imcDVepcwdd9qHLwm4L/Dlv3scVUVgvl6Zy2pgJwSXtoRNaqKVhhh6z/E3OsOAwXErufM54CGA3
5KEHz47c/a+jIdfHR6VK6vwSRS7VTU7Fa9XpVd63BOiTta54rqwYLzTITzQBbZtIK2p/UflCQ7R2
lSquYEW6uKgdPvhAgT0L8JOEOAxpJzfXyUaU2FXIubwsTf/dL5Awgjct4IoFmiZor95mV1iS8cM9
V88GEI3avb7q+AhWS/e/x/SgzK+q9qcAZXaA5/3fU8by4SXDzmMb9aLnC3ToYLqajIybij8Gx5kK
Q9ZSQY3HcM1kfqPQVfLD6y464lOZBd7u9pwj3TY9Lqr1OCgr9B2E7tspWjD5U+Qa6Zp20AHCRmZQ
FRo04fntVvF3lfix4YT3B7zi8/7nn+SkKK92o6vpWIrrceq4axjzalpRYGxwIN0clpHh0J6JfZy4
EsbLcAin7nFW7xTjK4dxUcaZS9AIGN1GsL+lXYkocfV3Bt/DMWWZ/n08ejbbeGkGlPgdhGv9s24Q
Cy5azXeYZajCxLDi/Ivh4BUUc+0+gLiIfGJcmNMvFd+ur4zpe2L+YDdcJoeWs/FJdzxgalr9aklZ
Z3yuXWQWAbGxThKoRNbUBMnMacAO3cSP1k3B9hhbIyVnivIJKnvHda6KwMktuyELHE+jFvm1NW6O
a3YekT3vHPj7h55sXeucpbOgctB0j8/jhy0X5fPYlA7J+X+AJgpr4a3UA7Mjo62aFxK9OUnpHT1X
TiKVmpuhKlA5Qf90dD5niiFH/hy018YfRSpjWO21zcTLRFNR527PjvlKIMTMDNgUJssDJ85M570u
zRclsZeVlhof52zX9O67mwF+VVXI9c+MYEb4BiwkZqp4V4oRUdqPrvPVXNZ2k4sh5sjgXrcBn2kE
Gnf7Q7stH1TzpOzOgqm9a/9ySA3OoNMZslVTXsuJ/8bQY0pzSmifSPEQHhEc5TirSU1vNZu1rkYw
wPrdG8EKK3xfEMFHZOEWCa4UvF4uvhdTJ/LHvRhqWBCmiylXSy1tFBxn2qU3Rexz+6xHovuM5tdo
qKp2HCsALgSrS12vFtojWt4k1xFLcytqNf++hQ84ePEe4mPwehXQid+JM0fEhFY7Q0ZL6MWu6c34
QWx5PWahic0IZxm1wRq2ntdxSWudZGKnBWVXbWgsS4drW0y03NBBxJ7AmuAXkf2VuLCV74/rD2TW
nS69AtmOPE74ImRWGXuu9AkzhkjE7iWsnEhdMBbnRmGqCQKQTYRUJA0cho6Vjmb1E56RvqMPNAqi
jg4ByRRISiSgWNWZBaOMPmrwYzyhHUJI/z9C0A/FPyVh3STRYfyeHElkAOlwUaSdaDoFe8DeAdIg
FK2wQOqhN5ZyiMw0OmaNIvR9ySNp9g45dEHSNVZvGwYROIwHLqKz+DqH+ZFxg7WPxykWPNVmemzk
lboZUm3CsvKfVrt6gvK248F2MEKCTVR/vUg8LGya1Ux9jxvDk61AHTd8P0VDh2EDB8+iaZGJmeUM
EojK3zGz/vLr9I5FAxNt/coIsxPYhKKwVUeMsMX+JD4IJSZQPQUZs7GSj8astBs7pN0YqC0m48ty
r/9mqJP1NFmV7Q2phuJV0V3Wa0JHQQxtEYNbCXCbb6VNAlstyr1GxRcMIYlvl52/X/e8OxV5VKfK
kBBfIBQdAqH//zWxhjYYZMWMCzMenq69OGMCZWUkOmnDU1iJMc3g5McgVOFHjkv+3cNyP7ztFAOn
VWd73otIFN3FGBErR/2YfC9EhAFOMfq8Oagr/Y/FdacJ97zE3qm/mfrC0UD+fE9ch8opZrsoQPBB
fRWsmRwh/Ifk/zEz1a1Hg+0qCC5BS8GeDnwsvNHUHsPMnSP3bl5kF4+WIKMCEUdqRA53OTBEDgNP
bKyJ6LOrm+uDRPG+kG4s0LrVn3ougVT0U7c4wMJKQfAG65xpkhOMD81AxnwSG8smL/FbMlfNa9N2
cRvQSCRJJIj1Iv5C7HHll9eJHAQO9tbLi9Ow5+Y2q/6EERZR6HD4IHRp5cvsHXWYgkvT64r14hYX
L8jGndTxx/t8Ug+ucyM+Ny5jPPJ834qX0zG9WUA2u3YaqZ+qSj9reQhsZwgsatktDSpCAwO5HrhJ
5Y7THwdofP/mGl4Al0oqFsuvaZ+02xIT7ivZBIGDelwg8HN5vq/oeeVHZ9fvcyAWZBzar/0D2Qth
ZWpTIGnuRpI9IthGQKZyNOxmtEG+CteWLz29ZHI6l+qlPhezJVFjIWfLAvmQy76YDtPVJ8LX8ql+
XPkHoaka9yylo1e2cYfCHEVZaELDAyuwAPtbg7ir43GS5gVNGvQEkClqx9rQihQY7XqgWfPSDklG
sml1gJuNApE+4o9yQab5zHxGniFFCjZBHLRrdZy4GShWIShMq/WzJXdgAswb2PTL12XtmAClYHOz
pRVgsST8Za4NctDV61ZMUhHLoE2p04mlGAClGHmbiC9GwwK/dtxlMZnvqVZEPbjOx1JgovJpnf69
IgoTTuGl+h0MfvdeMg6CZFGE2Ra+TNyuAWZlDg4Bt5PpFA9f8CZWAuSg2XuRLWvcmtRLW8MWMk0/
D0mqT603tAuM/LLMoDp9KX0u85PmpmQFp1T98EWGU4mI6lA0/K2qp8TeNU4Vf/o+kyxdTWv6Kkjo
FYg7MGZNJSOOxnAp79ZtgArdrzkCt26ofQgREogfjD6X8qOXyb+0LIAefL13xS00ewjQWrNaSN/J
NFUnAme+JmjEH8y1rVr04Q7WHwa+AISHoG97I6aPd58ZeQnFZ+s3AtRvHcv/A9VlBKJYKTESOTfv
lPguZjr31ZMwo2tHPv8HgYTyTs8uWzFvekJl9yPF/3W+Y4itAYXjlCuxAksnnE+EEOkNVntg7Wyg
oOB9LSS2/USAawuGdkpUewcbPaieRcRhtnBmmBCSUbTvRzRiYxTWRdmG5f2gig52FBhJwhOSOx6y
ED8kU085mMYIJhy7SgNdqWwaCbEBr880MRHVcP053yTNZtN5tZm198gCJTmhD35SJhlw8NZltxnP
zV9N6lmZPzWCQiq/7ys2qaZ1QOUMbS5L9VAZRVvT4pp3/wssq5XWTl3hA1l4AmKypmmHaHWUcatY
RzHxfA8nKA8SpIvmKhYYBelBhQxdnrJ7NQx61iG96tAxm3KwqMSIwXVI/H1kzbRhK8KELHMxLMZY
lPlaKHTV0pJpEi7RFjUhoAzp9VahmTgY5RW8Db4Eo08fimbkEQIsYX3CHKDZ2h60aJiwv9Z3reVr
shdXMhbqOZLNdbDZUGmzdS0mvMFHQgIzNPYH2r4sbLy3jCU2MI9vTp9rMjEjZXOc/RBHabrCyD2I
jky8FlPSdIy2dyGNttVKJmBwUFyKS9oyBLTN5d7h6DllB9kZoLcz8CIouyeSN8xXm5C3wmQu9RBL
rtovja1qcSBfmcMXQGhwG6ULTwq7Bva3/fl2A4VRh05vljTUi9GutUDPQd93kgkIIt06aWrQWwdC
z9oATPjVCp6Y1I6luImPrDYhB5e3//i+hVe4LkPTrxS9UbcTOZR6jrE0N4PhcbN3aseQo9SEpDEI
hJI9vIrows5lYJyxPVC6ZQGk2HtXaf2ac5orEfugDXAA9bZA2VJ7xK4o8TDLBzhLKhkFTmy7EFd/
gw3CKmVFh8aT1PbFpvPiLGWitkQt7W3wBaJopMKWibSQgmiXnk39W1S/7IvL0c9Qimve/wom5ToX
lBhJ6Bb8PydA8ttL6cu7e1m8xT/jBX+YKiOacq7yFefgaU6A09SeEO2Ix+syUaRBYrb9q1QPvHVy
0Vt+wpk57yUOu7XvqTEeiJq+WzgDzsmt6iRaWuB/Nv6QPCaxor10JNA/XzSGWGO4XIzjr3HO6HOp
gUErbPpzhRUr5u0kzXNirhg2tBEVbyLd213M0uas9PhseEQIEHgA/XTXoYERJggUuDiFtk/Hr2NQ
IFbOs701ZjWyRj1K+nCTAUB+DrMiXq8OuimoTb7BUs7xK8X8xiOkI32bc5K9cWKvH0L+luiVqZu4
6TJiJcCw9qVVYE2CztpN5iYgxI7nGkTRWZWpfTboZSbCNS+5k6IWAyd6FMoqZr/TFlpmzj3mD8GY
dzacb6kdrdenUVcel/gL6n8WVpnHHCZfKCbkWKd6u0gunHOi/Q3LHD629mr/naxvEsxzxbzngfUb
xWEBBniZlF1eYkFHm+MDB8PWmVatavtMSOiIYD/7yjK3UVOiLbpWrq+nAv2hWJ6KqX4IoRokBZSY
6eqRG+HTva0LvsXqS7QzT9SDxlUIPfd1i/QUune2Zq8qAeuweJ7CWg4bzHa/SzkncOhFgAlywFv8
Xd8+wmSet5wGB/yEJSJ8CKiiArHukgRupm56FsTpy/e3t0fBGKhmgCk1VPsxvRlTcGmjP8ioqqwB
/vZ2B2ByBUMzL2hAm+CJjmtFGlnKoKQIEDTjnRC/ecsPjgPrD8YNogQBeiOumk9UmIVtJatHkLsN
peM0XVofHV+yw22Op0S5xM7U029CkPQ7EAlPrrZ7Es0aoU7XRRgBZVD+F8bdeWiSkljm0PrqtjJX
ed8/EMtP+0cOe+nJ+oqRt1jcP60OaCfolOsDcfrFoAncmvf36wIlpKbpx9Mm8IQE3n3Zsmc5Jvt8
e6PPK03mBNe3Mf9DyZkBHfEPznZ1+ghxRSWerSKGAfPMKZmp3v/xCmQLgAsy5PUo+3IcirTTGnqg
vZ2h4pPf3g85R+Bvc5QN0qNuQRiEiE4myEa+0AvdVBaOC99tGD6K6kGslhFTFUWzadQiVdUu/z26
KL9SUHHbai7JNa6DamL0eCAv3O2NxrM/nLTQLgB5H5xOOHQJt8IhgJ6XtRuMwlbVRPQFIQRw1q1m
9nGg62vrAjCAuTSWxkRg3RRg+fLJauTK/A2nC/fUNkPZph6l146NSVct/jlMs8FG3TumzZN36gym
xTe+4WSZ4hE4w67pQQfwst7+S0enAdeToeV28dFjkhGUDuiDZmmeyZyo/RyZ7+2EVhaAPmzk56rQ
diDoQd9hKiJfE36CP2TiefuYn6/soU9HeUmfHE6U9Jf+MNujFzKr+xo3JH+T9holajXNv+XHaDUi
6HejGSLbHAsTnImAZgV+JTSHoKzx7zilRZTihuaNL3h7cXga1N2HRTClfI6FgVFANlSDfOZIKCIg
4iyr4tHn4RmRo6oQ6dizhSneNWR0qDZGrd2aAnYWUeqr0UxrvH9wAqeEc3ZCCmRaz8sk2O/sYKy8
RsnYRUPSmgxJ9r1jKGKO/QYDTpwkOTNi0KbiCmvL5uBiloIToVFpz8k37hmT2nMYGJg61IDQjMM8
8MoQFQiat7G3bJQPmmgOs/uS0OSNYA5CrAMmvmKYJhxjETyusYal/mjxnpCKo6/FhTNq/MBe0xMx
XDgrOxYLUzO2psrxz+RcQY9hvu+v5yNNj+uY+BIISq1KkPEDNlJkumK+mt//6Rx6y+j4GmU1Hzhh
ZXnIFqA32YCXUPxhQwlaV5ajQI/LI+y1HDIwSn8Hq16VzE4GPkaJynjfnEJGndeoezwmzoHZtoEK
k6Pw0rQZ7IY0YM5LrqA2104pwF6FRH3odtiWCfPHzrydo4zff3N2aBpbQ8V8gnX46lPY+0TQR4Ej
Yu4U6l4OlVpbQkdDOif32rSM/gjD9yYY572wIsnyIh/pQt17tObYZ1pSX4wmqje2WTaM4/oqj372
rqsGS4wfdFm+oxXkFZaI//YRQ8gDSxAj/vq7TA3nO1Xp5kjMABV0nNz4i++J1RfxrKg4pKm3J8ze
M+9QHeeOpgQ1qJnK9HFUEXha37+YGpHxTrEurHs0tWg4oaKenKucUuPRpMxCPtjQamckjn2gXHmK
Jj2oDHs5BWOTtidktILgC/kZ/zKpLtu1S3EXSXwiZwwsxeOZetmkLvmc5tY9K1dX2R7i/N3j/hef
h2hJNpcrAIPYxxTSqGrd8tXg0YkWbrAKmyJbeMdOYzR6Z2q5urMZ7IJ03XgrzdvScu4EYAM6b1e+
LUPzII5ZqRLUKjtwIXQ/rBdUBnhULXcnzBMPrWzDY6MOwBPkAhDB6qLJYReOvJRACSPZnrD0GKhM
PkwK5URV16bTEmU4/O425TEMed6/qaAKIdn2DSrOXBHsGRMEmWVH6RQpddLjMu4r3xe9z6CgL+Su
jgAmM+nYGcBIeF6u3g0b1DsIxk5PIdrC6wePexXIj5HUaPShedEuyPjiHj3qK+RxBQ7kcYr3RDWX
MsQ3UlP1t53BL1ZKcFc7emk4xhP5lVCLOBg3HArcIjYy8cMylcpsOXByXig8Ak5FZMnQgX+p6rd1
/kayBZETa7KYbh+0vTvQpD1V1S2twVnVYdY6p/Bm/KnZCXdD/Vas6rraEcrVSFLR5/jjJ/V8DWXJ
5zTfQI/z0uiZTIO/5ouqI9Fx7mkXweBUalj0U6J4nEjT5Bxy72ecXLzUKixv0/8jwWgzUQ+4Zf78
YcwNzjkCzSjFXl7qeTRCGq98OPZOmjFBn+ZbjQ87G39NzUogB6SSjU3VYv544Cusrx6IcHjRZgsy
hfRHBRCn2/65Ozcl15xk9x7mIpi6vkDiOKimo0Nv7d0efFeXUbhWRYBQFC2baIDfmfJEiNmPPI4n
sOyK8LALsRY4+hHo/iDCaXMC4TCkC/sgo8MIbcyUU9jJ64Qx9QJC6icjsmMtRw8WRcfAuwgBOjMQ
kxYVHU8wpbDo4SWOJWnP2w8zBR7UWiAVfJz5D+CocILV8iEZEJDrhQEzJKIXgh21Mompn76FyF7O
FRJy+gHBlMMlBYgm0nf1pKmKkH+TQbZOMI9IglwLNmVnAwPi5zXFPPJEZXP7XKeCDLB4m19ANrRP
MdWczCO0d8Utduj3lD60gzZKzJPsdg9DakrYo/Eq2WXYAkxO/w997IytJqt/GRxNgjRCK/20sb5D
1qce61wi2qQRQXmeWcXVRPK7+8y3Q3SDj+gqda56Eb2P0zjM1Ju997X/WVCMY+i9tCIho32mgHuv
X+J6BqITqC6bFps0LrXlIm/cu3gj5PO5lhJtSOzbboN7hrUMCwOaz0hyZvYG3FRkkAiQ2mk1wFMv
B/Su6eCs4DSYS47fvbhwvmMWgq0rUXSxzldoteToNh+NYwNUqk8VWY68uSjIdrAYWVrHP2QI4E8U
yD+bEAonshhQJbzA+/VThxjusPfoQOJartEjd6A6jP1ZBHKorbOHfcAomMxnVKFZFFnC7NN9OIMi
AnQ/JblA6AnmUMTVW3P8gWxth2kMGFkDBkp4sYcGlAX/OYMnqXkGDigr7FR26N7e0S1szZnjkbLO
saEop5cRxRnilj0ZeUt/XkTzKJYDKKB8hNCHV27V1mJqHWJrzQSoc8cSEn8m1KtJRfKl75b1S3rS
tV3N1JjREt8YSdplxuat5p8Y+ySTMYa1m1o1cCFKwf59YTd4BuzniFERhsnU1hAFg++hqsFbMRw8
aZ0O6GIEMmmwIqAnsQYLqV17daNNfzuEXfP1beHwj8GzOo/ZaCNPIrD8pirp+a83P5ueWNlzvqRK
p6ctp+xmpLrQHDe0Os/exn2Myo59N+9C+h7EqpR86+42JijhYcoqEcBhsCkcaRC7rQf7a/hFeCLh
7c6y6e5cEfqt0t4/7Cm1MvB7Y5+WATvj76bfeyMa5pNZyxkjBW3ADl9lQ6DebGU6ZCmT8v+u1+Ih
AUjxU7J97pNwQ6FxJFnGHLQqHDCtJV4eVTgRhMmznGWQh3VpWezeFTORhlH0xU4K/evRrQlMhr28
zPcTZ1RZDY2PZqCfA5BDdSOCVGbpwlBAFTYRnf5M8cHiFo7vk8aEN+CrUOj+AWp8BX152ufOiC43
8s58+g6z0USXmFVBjdwZwQ6PDjg4IJuSy/AVEz9JuUuloEEXHxEfRzdJJEMdTQkCiD6QlCEVsTtS
qg3gc0criFWwDOIUtOKyofH4wOzM1ZLCm+qJHBNLyFabS5T6dtLHuTxARS45H/Bd1wiU1TnpM2cN
Oz1MwslCQ+qrqptHrkglWc+8jgpTWUrNsATVn9eJksDK5BqWzNUQEZNpNRr3o1nzdXd2KFUDNXBw
RPumqZRpFd0kIxJ96QUgnb1tLQnTfpDe2iSF82nMP4xkjSfXQhwMM+WEU5fgUDYoego0vusMpJRt
MZNzaVaOsLu5AvSYrduJYLnrNQ0UV12oAyEc/Gt8GM+4qmYNqeLcsMTUsjKDStifqjspryzimu6F
rkAqbivhuzn3xYar6ssWatU2ph9torBKMzIfbo+NmQREPFKvx1N2KvKtbRUXTPqLzsL4yot2VFAQ
I+0rNNEwNemWgZRGSlNT3BJoTi88AuqFPveQdPIOmV844slny9AE9dsQV9w+UIcR7SMQSPaq3Zri
XOVgRcQSzwyAiE80+HwAlGY9MW1OZcwon0iwSsQUCgPqknxugdAbqgmuJo5EKl1/NroNWTFtlPhq
htUSvtBbohQ1R4EDMSSO9bZZsNkPz5ME8MBTztMuNwS25QKrQnPeIX6z0Vj2C+Qxu5UOOa5XDpRU
iy07rbstiCtlxsd/Ju54dlX8cOhwrAkk8j9T/OkhUM1M7cykohXYwEoFOVEC/vrYlevzDfFUKSzL
GTWj7QumWKNC/tQG8/d3/vpZOBnJD5aks/oFkSt5F2xamcxcv7b4ABoyziXRA2IWG3CrdsqtvcGo
feaC8KIEFxhSGAwj3cV2eimCGj9cMgIuqZnnZprddeVfI6W8OYZwef0rhpSYpVXqzwS3pNOt+Up4
U7jrWO1okWqifCeeOp1Otee9ri1ogjQXubqqEsi5JcX8xm3znynlgND1PskNnI3XEosP0a2RpDuz
8mmUsKD2DLLNMv3Z7v5NZAq+J525Gkh1V5w9wzx0KUC+8hvXMtcWmA86unCHbWuJaUYmlZTIM2x7
BHjn/bNR4mMG0EAOBuoLG/Q0Xp8byhHAKm6kUrhHuVoNpPjTE/Y67rrxQCIozH6BdmjrOqUJD8PZ
8sozAI5yi2zUt1GTdWN2IxDokXSmLVosubwo88/DHlJ53Iun/XGJfznvI9ctMzLmOcx9Xc9aewus
XewXNGdH8DuRL/StA0jGP68bswyaN1LGvRA6NMKA5CZDi+DmAMS0Bp5tib5oGPwnszK+Vn2656VU
KA8b0sqEyaxqVb21WGsUMfPQ7lQDDh2r1PTkcZxhuWUBcye4xIepnIiwrElnR2ghy5eKP7lI11Jh
DdhHqWGMi/RkLR0m2eveC1IF7mya2ssnj8ZO4PiPo9dXWg6V6t7x8VprRhH8Cn1ROpJgjdgvxi4b
S8tTvEXlSXdfRkaNxbBEVXWWHCHxdQ1aWsrW+Vv4J3kiE0N0+EJxtDRF0Sh7iS2P4LSvbrvT52xB
1U8KkiPeBYgPtOV6CJIvdw0r9W4gJCD9H4BD+5gXRgMqXWWRteHDA3x5WyqKV+9sxkZzqBVqsrjy
yp7IO4J8xJvSnNiv1eGS4GnqWqHEMi5iShdVlTyEfr95PKhCkYRWKYRc7f0612ENB9ObJwKFB/Vq
D7iXm3cZKV5qjEj88ynopSEqvJFeDqwBzyMgpRGsqRnwTT2CnHtEzlLbcpcUgp7nr4KJBykA10pL
ysnJCAaWJSF7HR0VfiLbX6gTLmHO0nQN8Tv9RaAbaJO8h+0NIoEBmwHkk6BaDAY7XlK1ovZDK+bl
a5U8QCEArl6+0O9gffY3g/hBYkeO1+jER2fy9W3xJpqdOI0NNqXVlLj7AT8Paz05Pxc6+T5lPjMy
/TlLuW3oGbtQZEoF1UzYLA8uef4vap5RgCXhBDczZNU5aIY6HDI5Uu5PFlN2f0ROZqD9ueM9F/0x
tmZc4l1wsJZ6sZ4X2e1UPsitn2bYskf+52UH3cL3jp7i/hDgkERG3MquPCn2/9DiVZ+NLPAT35Jp
muCXl5KVZIHQDQzhiXXczL77HBIs7rWH90iTWhDvDv0xgtFiXTV8j0O9CJx7wd06FboFkiYzehWa
iWpnqz1+l3P08vyGf10cIWIoL3QGoCaovdCc/W1v6ZPstAscuVjK8Uu6HzOcJ9KxGpHfzuMaGilQ
37OEZuU2JT37fMmXDDlSYsNq3oRHZckcHeLbl++1J/I/8Olvj+Jn4zlq/kgxeP/b0XpJd/aCNAAh
M5cNIggA3LagHe644L12ozmPYIK1Bv3u7cJcbLKdC9EZ3Pfw1FPtnzPW7XYc5MQxP4rSIAa02jQv
mHw8HUmGXNKeS4sjXWb4NX+qISZtBV/KB2o5ekewY8/XtSBvjJ/GMjEkpxR1sEwAga+y7EE5YK2C
mgAX+KMX6mZLmOACUpyADgAj5JZAtKJleRxn2bhzepYZh0YsHnTpgOeJC3YafhOVULVe9T1bBZKw
eFsXovuGnvPbhdhCBcK2pduPtQfNDCHMwtx93bg4GrjWAZ7WriXCgMbDxSj8M66qEAgKUyCdupeX
F+qh0BbzQJDPOQ0t4B70wzcZ2S8xGv4OsYzuQPP7o8Gcl1aeDWLMnXBhoNz1IP/Elg3fSZ3QstC+
Y4NWE9rDq/0PFuHCsq5kDPrFqEz1qHLBaKvZSJg/9dVGTrhDgmeRbk+N5zN0Cr9NomkrY9ELrkr6
8g+GpFqXzvZG6rUfIKLcPC/5XTTiuHJIXMIuTBpCUrUQDsQU+vOqIWepv5+KKcIpq7QT1a9Ut+hU
VVmljXAiZrtRqOKjo7iM9KgeIpRc8OshPWxYcntzLQfIHiiZhunVezgX7+gNTi15mfazbsvCDbD6
82wKAHLc8LARMUMDaj9dXMBQsNYyd6rEjzZmMal9tvRITAxcr/bTKqNJYrjPwgQ/qjebNqrxlVwm
9u7u0qWzFCfTg5ww5vwv4+8EKdU6BebBPJelWp/yCPZuYAqOWjHcpF5Mc0zSDSrHCDuT+f8R2mMU
Njm3X7rvX2SxYGk7mgk2jBBOIQc/j9PLiB+6SPXEI3y+4PX4ZUK+Qkofs1ek5irhzUZU/wFX29wF
y4NL67v3HqYq3hVLO5buovOVxLvvd6TwSyunhNHDeHc0gToBIO+31JmX144PMNZVlat5Do9H7AWZ
MzTKr10xzHJiR4W2wPgBa5hqhcdIcKUB0P09f9fvcHjq4Ul/oFyrlUrHCRUQIbnmGOJKyLHkgVTj
Fg2bZ3ctHiTqm0efcD5PEnTb1Ksl0+j3Ki6BjWTaDR+Rjp+g4cXwd/+EusAg0X+goGJr6aJn2jaO
KfTdPHh6djnJMfJTfXSEpJfZxarSoyyHoy4McflZbWpgKqOwq4Vx5BgtY21YIFxaV894dk/n7Fvh
3MrlTSg6urV/iL5v4sUIu48VbToBIrfY+kI1+JkDjNQXUm5zOZ5dnoXs4Qrc33bFxw/TTOB6P0BL
/EmC2T0g6bvvLIYpA1cb9qVlM1+rtMevoY+FKLx4CEvMaTdt3WT0UC7Nd78yDUuHzWHuKlzcNpKu
OM+eix3jnUADkeKkMTSs3aYFomv1I/blATfde9P7MT4vxLn8w7JsnXT7jAibLt3Jvv+o3yD/RPHJ
fElWbbSGuOhgxrQ80s1ujzqSSU8TH3IpyiDNpiu7VWtQv91DhPEHFtZq0nTWe3JS+HX4p8K/aEnf
2g0YFdWiMfJTbuMan/4p8GoIF3Ww70Ut55OW0m54CPJu0tquPNIIbo+UPaxzpRDdiGGLHjkzeGdQ
cWmqOspYSbYTnDznnpaWa68WK4l23qIwcStIRxZnN46g8FuRbkG43FW0xiNOaYYqSxhl8kYESZK7
zjnFZRPqZGT5pD/Q89unLB3TpeEaNqbA/AyP5wGHY/fzNXXuoLrYaFmIh0vZGfBtar3lpcv85/OP
c1AGKwl/c1oF/B8/MvNQ68+60dmhwC6xywYHffdm0xDu3n05ayEhncN2/q6PEgP9V+QPhG8LB/Ay
rTYwvj2n6i5HhNoR9DCtzvXfqSlo10LCq+JNg9tKWhL2bp4YRr+jL1ASu7EvfFNCknBCuHvKBPyV
IJ+BuUSVM96D2sK5k3VN4gwyIVXCdnHZasL1f+t48Jouh1rEBugodaqQ6yszWYnRAtCgJkzORrzs
UMh07po07gg2JuViudKE+nSZH1OGCCXY1qwwbka99YSjvV/5iyf+5EFYR5JkM7upGo970WeaIp9C
IcDDcoTR4poZ2V6Ze5ay/dLLMrhqHRqnG0wOCk2VgjgP89WaXLVA4TFoe1fwyG0mexMy54OtmkUr
o6xnzWGl+TPEi5mIuu7UaJUaM84KZZSa5OhRWR8sLTinhFNGLKxIZ+3YtcJFQkUVupF+accbmL/O
PXwctI2jIeCIpP9YuvwksAHknaAPvuNsj/5+dnNFgdEyB/EwCF/Qz8Rylkub0c3SxSiJ7IX88/D3
4vcFOCjLOs6GWHQGYqpo6mqqPWuNb+XFYBdwx19fnwj08E5+sJEj7BrMEX9ZYhUjvD9n0XD+MX1w
8Ba1+938usYu5+4MktmjS34CFIHw91YADSQpECyfOyNdAdNokyQmUZnrk1pm68lLtBbKCVoXlK5T
Cf0fVvegW17OQ+zzb5iKtzWQT5H+sT5msxOg2SDs4nNAak0plqtF3z7YEHqp4YjoMssZV7DV1gHY
iDGx5iCL6mSatx1wjkNQ1Ru90l3nuhmWk62vXyAho/eFHNYm/vVYRn6u7EFERnQLqQ+OWzmtRj2V
pvrnJEtlV+7AT8UZD9j9FaDo/FdSkqXeChp/9nL/0mi5vgd4cBEs9KRHQEbElollQVuaunaGJ6/D
XJ+aNZ/PB6eCjBWuMbOA47UjJBuMuA3u7Fee904sE0TkDEmD91FuaEY+0cpjLuH/nMhqccX9EwCE
4owNn3D8drJyoL39yxmoeH59PNdhtWauG2rCDmi5n5mJtbTrp1ksJJUhTuDOh/IJef6oMF+hHEXs
v496yDlrbjYtUIhM3LEzJhEwXen8v7zvZUkhv4BaqbFcuvyeaKDuCwXTsF4Cs2Nn1WgBfjC1/cPk
HMBvCjHnS0AaCjaZB85KN5tjN1YSqwFOoLqSeSE0X0KwiCg9IUQ5sTYeJYN4bbYc+vd3PYrbQ6tN
7xe7PARO+GhZVEUb9URCxYH1Bbdc+FY2icx40YCFiHdvzDZwwGfUc4qWfX7rbP+Hlzw6+iJf8UEr
RzQ5cLgJ39EYjZdIoAYUC0BdSVfebZL3HaUFA8sG5ZC/pbi4AWaHo40ZybF2tx+bmNx/KcIe5S0t
SBMn+CUMXxVImcvXBcvTkV8COjix3ajuKdlG83b4HBURus8bX62f7cwCepuvVjiabubxgzhviTYL
JsueC02/38rk2NzWMN881hd9ilm5NXDUDgbzS/H50A05EhkCFXijQL4PYB2BM6x5Adb/9wE5DYFM
TRw9fdEPT6FWxdyQiIcRQJGxvO8mO9Tyn5H1+HokN2eoNOMFBWDjRUYcgMKWyVlkI8xgjtgFr0/J
5pPws5LDv/JbgeQ3oReLnvacXM5iJ7g+XJ3tjYZCTo5UPHrgDHJ28KcvrNJVzQeWn4mFDb8Rs0em
euyh/jM2NSctk5BkBHqsM5J6n2OKw2TVCZ4rj9/2CTUrMOmb8W/TZBDuzdW4KkFr+RnO17kanClk
toEs5vwmbPRh3cqC/JnlQyqe74/H8D/K1F4oc42VdmwVRq4dqMyDrBOv31j2ZYwew13ym98wPzWJ
5+eykv7vHE1Cz0aqlvXucdwcHaCJXXlqJzGqdIEKvlFYAKssq8cHXXjReGuYGxfva5yOPhwVl3yB
3yRfMhH9g46D//pow3rBsLratCip8B7eayniwKYezz/AzNZexpbD5wbzM4FagNiSE+trzE/9KwQq
Ri+ATptNUOpcEuTQiPJ7l8ISYNby1Ad5IfN9OvTmTBblBKP0Hj1Q/+I9Rz/0J5B5+h3L8rA9w2e+
P+QGAqoUm9vAjxTJbPGqxsARMYmgqnvjP1TCpFwgNPBqPBFPoBnQXod6u5WJKIwZYlMULsLZ07Jx
p72vzXZ4vKZJmPGzF58cywO/Ba9bsTMTUCh4wwlWbHRroj9y2dw+Hfw+8yGpE87CjEhILxw+UHD6
lzHKNO7FihekzWn6xbYglOfyK2KQvZev2TTOlB1NhQmFm5qORZpCRRusZLzaW6yNu373iU4n3KH7
Wd1v63tRrAV8atDa9qLnBykQDJDZVtCsMcqk65FDUElizuynZ+YpXnpv1QLESOcQnoZBtxeA06GY
TaXy0lILUtdF3015HUcZqKa0ps9A4E4WIeic+wEqaLfTUia+ULLjzm9VVd/1h7dhXXqLmaMowh+B
YgE5Mc4XLmidmsxa3aDGQrzK8nwYTZg9ocwxLxfSDnjt3z+aoFIJaAYBbGXAhRcJZYnOq6zJ2hPK
6UhfwwxgCz6gGEpp/kBwvXLQa53aGNqXZ+7pLuzx1iCgzINsuaYz2Ycnu9X7Tb1vyZuo1gO4u6Df
vBxt/e9Dpkg4UyjN3r4gz/lL186M2rhGUCNS9gIGRklryFIwKH5FgJVUeT/YS6SNJ6kTD7wcPki8
ZuXcK9co2p4CjTBRRadEjG+liqxY+MpyFkhMb+bGrdWgINpdrR8wxrJz1UUNyba+0jO2vxNw2pi7
+yTGeDztuPapz4/YnIrZkpH8L6YHLjkB+BVNWMwjRXZUJHenL7bFjT4dauNCPerOWrvyilGI35p9
YjbY+rrLz4zQIDIs8MZLEBe2ILgxdCXbKsAsznzx5tz8wV/OEvwpQwyD/Xx9IpDZ20GSkPd8WUcF
uNRAxTOtkBii6YJnqJ7trWyChIcczlVDJnHq68nuXvjQP96nIMmrTOXMjGkVb/R3gjn8ir5u3tzk
F5aehjgko1dgVakgq8Pp+JWkJadyPhQ9KaMgfbo+jUl59paHvIjpBSL8iIFNxqr4igECHIASNeLq
8pOgWxRtVVHwUBYMrL6Q+lM+QBX71mBxM2MaG1sNCMSZXRoV8emAxNWAsbC7xKeUkHvKJjNE4tyg
bYMZ8t3Pc4zuQWrYwbyEMS28oEj28hEJzWPhwbyzp6QuLSFdg0V/tQgtFKQTZfoLKcGZDW2g3c2+
Wh/2z9LympXEMNpKcvnYYltpjmMNIw6y0JVmSsxvojOJGnPQrdOS1ANvRyyJf1DcMALjNsx9QQpp
MD6LoJNAUUpBOROOGCmhHLXTrGVsu6JP6Eq2nVjkwPIGbVdAtVuJO0n4pQaMZoK3hvMpbJYVeZz4
xQRtw8UUD/IZOzHnh/4NUlnsxjWl8aUo2oum8Uu3JzaGF1I/yIItfsv08QbiciSy9IhPh04LWzAT
5b8uj9SSMcwOm2pHWt0T9xBICxYwgfnxbGPgk+0O6wnKD9WnT+8QSse62mkOXDezk9ts/kPDWLl6
YQu83xoTent5Wa9QUiLHPkUOnLaXuclYYQaP8hFXSmhG4yvzv36ayYHPF7f1Oy06IRK8TFvp4Buz
ssHP2Qm2v8sV5PiKrqe+7G9q5e2BcGTQ7zbLo8cRIbTxJBQjGKdSOYTqMItePzZY5bMh9SWgHSeW
KPyJifArOsxW25H1/sVxGaczp1ZWM/5HfkU08pclWFRpG1F+FG2lkdjOtDvTMhWvsfL5A2DJlsV5
QkQQdGyb9tUF0emFf5EunzWANnkHOqno30ZEhZ0/AVdnuhY8algrrSwN51alyE8Wm6j5YPpb820O
eV2Env5k8eOa7irjjrCxFduWuA7kfAzPtJTFwFyiYzPZ8lxJksIRun5UWkV236hcL9vpkSeifjnX
1UNVkewMz9oQAWKsl1OOJOKMEk0xrcmk2NF7ldnyU9yk1WZuf03SlpK9cQCyoMvDPY5brqNOR+Ym
0DYOkyVA3MH27pYxdAyZs89CSxuPLF1NzELa497dIFEaNjmFDngMmZcmODDwy22AfY52wOwA0CKi
+DU16rOAakpBEfDtXmsIYclYqAxhN0K7waWWPgdFZ1bvZWMTYa8ka8Df5pBHiL3LS+UaNAMvDGfi
zQ==
`pragma protect end_protected
