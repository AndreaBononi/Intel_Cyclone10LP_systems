-- avs_hram_converter_TEST_basic_tb.vhd

-- Generated using ACDS version 22.1 917

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity avs_hram_converter_TEST_basic_tb is
end entity avs_hram_converter_TEST_basic_tb;

architecture rtl of avs_hram_converter_TEST_basic_tb is
	component avs_hram_converter_TEST_basic is
		port (
			avalon_slave_address         : in    std_logic_vector(31 downto 0) := (others => 'X'); -- address
			avalon_slave_read            : in    std_logic                     := 'X';             -- read
			avalon_slave_readdata        : out   std_logic_vector(15 downto 0);                    -- readdata
			avalon_slave_write           : in    std_logic                     := 'X';             -- write
			avalon_slave_writedata       : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avalon_slave_waitrequest     : out   std_logic;                                        -- waitrequest
			avalon_slave_readdatavalid   : out   std_logic;                                        -- readdatavalid
			avalon_slave_burstcount      : in    std_logic_vector(10 downto 0) := (others => 'X'); -- burstcount
			clk_clk                      : in    std_logic                     := 'X';             -- clk
			hyperbus_clock_outclk        : out   std_logic;                                        -- outclk
			hyperbus_master_chipselect   : out   std_logic;                                        -- chipselect
			hyperbus_master_data         : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			hyperbus_master_memory_reset : out   std_logic;                                        -- memory_reset
			hyperbus_master_strobe       : inout std_logic                     := 'X';             -- strobe
			reset_reset_n                : in    std_logic                     := 'X'              -- reset_n
		);
	end component avs_hram_converter_TEST_basic;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal avs_hram_converter_test_basic_inst_clk_bfm_clk_clk       : std_logic; -- avs_hram_converter_TEST_basic_inst_clk_bfm:clk -> [avs_hram_converter_TEST_basic_inst:clk_clk, avs_hram_converter_TEST_basic_inst_reset_bfm:clk]
	signal avs_hram_converter_test_basic_inst_reset_bfm_reset_reset : std_logic; -- avs_hram_converter_TEST_basic_inst_reset_bfm:reset -> avs_hram_converter_TEST_basic_inst:reset_reset_n

begin

	avs_hram_converter_test_basic_inst : component avs_hram_converter_TEST_basic
		port map (
			avalon_slave_address         => open,                                                     --    avalon_slave.address
			avalon_slave_read            => open,                                                     --                .read
			avalon_slave_readdata        => open,                                                     --                .readdata
			avalon_slave_write           => open,                                                     --                .write
			avalon_slave_writedata       => open,                                                     --                .writedata
			avalon_slave_waitrequest     => open,                                                     --                .waitrequest
			avalon_slave_readdatavalid   => open,                                                     --                .readdatavalid
			avalon_slave_burstcount      => open,                                                     --                .burstcount
			clk_clk                      => avs_hram_converter_test_basic_inst_clk_bfm_clk_clk,       --             clk.clk
			hyperbus_clock_outclk        => open,                                                     --  hyperbus_clock.outclk
			hyperbus_master_chipselect   => open,                                                     -- hyperbus_master.chipselect
			hyperbus_master_data         => open,                                                     --                .data
			hyperbus_master_memory_reset => open,                                                     --                .memory_reset
			hyperbus_master_strobe       => open,                                                     --                .strobe
			reset_reset_n                => avs_hram_converter_test_basic_inst_reset_bfm_reset_reset  --           reset.reset_n
		);

	avs_hram_converter_test_basic_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => avs_hram_converter_test_basic_inst_clk_bfm_clk_clk  -- clk.clk
		);

	avs_hram_converter_test_basic_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => avs_hram_converter_test_basic_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => avs_hram_converter_test_basic_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of avs_hram_converter_TEST_basic_tb
