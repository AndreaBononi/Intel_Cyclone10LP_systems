//__ACDS_USER_COMMENT__ (C) 2001-2023 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
//__ACDS_USER_COMMENT__ ACDS 22.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
BLMU+GqjlUMQQ/SWm20iPSV8dpIFK/qpG1PUUYxij5Kj3ypaetwCKC1jHawAMV1b
rMm+dz4xJfVO4xwDqFJSUSYmNrpCN5o5/yibneTbqA3ewohpjyETr9gMz+mHKQJy
5jnEmkaS13bUhqn2blEzM+BilI7K9120OkhdBwPOW8CR/Pf0nPPRug==
//pragma protect end_key_block
//pragma protect digest_block
JJN/lkn+Uh/GV5Xr8uNdYGrPSAs=
//pragma protect end_digest_block
//pragma protect data_block
UyKwxpK5HNAQbXCs43EUALiWiAzoWDX18/Q7LKlNKpyWaT2l12ogLq6kJ68U1m5n
ylcl3T856+bvb2umCoMbVpjVpw9Ndume2ddrdy8JavOt25E6Pz+gjCIJNBAmmqGC
StqHPJVyJ+jww2t46jpXIvpIbENtBQ5mBq3g7R76G2m+BF9oMmNO4IaCNE9XHoOz
eEn8R6CoIIikLTfVWHAmhJzl7gvppa22J9HVbGVcuEp1xPTT3/aA+ELpWv6CtEmI
81zdPo/ByeBQz98JVQAQnFL7UfEwAzMqFwwEbv0+MrIr2ZOiSy0M5mD3nsSJ/TO7
quzjSIEKWg0H4nRRPNdyCyErbHLwT8aGRbJ+J2FSKHZxEBe/sQf/qSQ8jgQmY4v9
6YqXhg8MGsrLfaobELa+QHqX1wgQj9L5fiu/SycYyZ2reWsL0Kejsjd7V3/5CaK+
77yx2eYYL/j4ar00o9muUc87LGqQgxJzQZp+xIPCVXL3rHYfAC39wUKwC2pmnbOx
U+xCm9EzB34SfJHKDI0oK05EbSTulIxnN2s5YrBb7ZXiDeLLqD15BdTi73OHpk4C
b803A26bPX1NRhQmfaYKL0W93vAm2WCOIifJj/iHUJtHDk+yjyEnejsOsvXNG0RE
qiyU5ML8/4X/Vogzu4GHVG+A5e6UxTWeONG4DPd+OZw+eks0qhhV4cXhxZ/MAqxR
sNlyFfsACV5RAoQwuRhMw+x/Q7m86VkzOb92fs1CwZcsd4kvxPQgghqcB4YIeITm
vixEwgVT5r4fFg7vF2CnAHYVul5BvINCPBISQ5Tt/VL7llmJ615cCWuju3DkEwvD
fArvklHugIleBouMyCe5n6YCZEmmImXk/tdyyk8rEavmeMUR//tJmas7I7Jx4Mgz
vDxSOLGchpZU50WYGPSbdON1/jKU5ikRO344OXuFtsQXAPd2mCvE5P8n3XC3Z3rG
H93GNgwqoawjYFNNCS+RmjFXEjPOvf7kdGp2G+qPXZ/VbS2JGW4OxlQ7W3lt38WH
Ba6/nuT/p70nyun7ZWc803164tjAPl79JFTPzsZCkBMwRpxK8nlnvmB69tDEm/5v
P9kS13yCQMes2hp50sQVuB2nmKLNeN5hGtqv1/tCboKio7f9ORSGWySYD/2qblNQ
flNZAwGb3SkuArT8THp+7oMT/yh2MJiEIK2AlZuYkKJoMgm2jf1hvEsVidpO+5FD
fRpdC5aflM16bjm/uGhuBV0xXQjWeo6ICyHxRR/J+hT3EhmcniaNsJSisx2mlMAm
Q2kfWGAqntqO6LwhTQkstYqezP6NNjCeRlWNttjTQMpQMp3FWfDhQM9KcCJgmd92
T6ehUXtgpi+AYXyQM/6/NIp6VPxB+Jc7Bj1DZWoYJ/I8l+zPP1QNknChgHuzKUg4
7m12fTtKB+h+wtosh9s6Fe4uMXtKkmZDcX+q/S22ySqiLcuxVo0teJCUDIXmB/tX
MI/rtI/qTPdQXSH2uOBR4FixRo9h0abvZ8sRzT3c2Z91FuyHucWutNN+NoLDT3/M
E+uO8LuBL4jSwiadccX2JKz3NvEWWHYdy2PR64yalywgNArcHlecsWoax5CuZCtk
Dei9amMfSWv+xFHqejPPp4fWpUzHpfVWUWVjb2yMsYeMT2Q45bOyhXngAAfQTDwa
V5Y53jjC5CVWWUOVrSf784zZ+FeIEzq9Gf7RightFgz4EX/vkbmA8FQQye2MjyqO
9gGjHTYoopcEeL4bHNC3OaTN3ryHcv05G1NxRNlPQMjCnWUtstCFuTppnmmVl5vL
CzIVvP6d1Rg5BL8OCBG1y0+EaAIa4RRdMpgUsZaCqH9K4ll9Irpu0OBlmpBXYT2c
G6A5yCkYEHCSe4z/dJim7//gqNc2fCW+fUL/WgT+HkrPb0xIOOrZn3W9pWikjUoO
LAQ1Wi9aQyaNupWLXX1ReMnxUwaYzZ0sidknrDqCcHbdbksY6SqJ7eLSYME5sADs
+An50Z+bX59+TdaJ0p5+uq6D+MTvib1lSV6+UnzsK3vHEI46ZzT95bGKGpffWtq3
CrxZXeh3YeTXBxE+0nXUOlGdjdvMY7vLdPA4NyDp0Dju2+QVpXKU7Aad8RzV2wQa
Q4CL0N87xeOhUrDqZXOJrJF7CvuQtxvFAxEQjRm37o97cxyYsxCtShl1rzqnTA1o
0u6iCNd/RT73dXSMIULbcWr4lc0/2ykIyClO48qOeBg7Ii/qGR9aK72hciG5t95T
G6BsYgOJJSWuzohX2NDggFTvMeBEdTfZs5pEg1glODcgYkTUpR29XfhQrDN1FqHZ
8q6y9sc3jy40QHuRdIBCwgfQsBuW1kSharmvYX/glLLkGSmmlht4aTIMpibLLMj3
XPDoJDCCSHBuh/ozdKbMeAby+Y3PHw7xDl1R+Cf7jlpb/xwmX9iQreQBeF+BPPaP
ghw0CEAjnyHo8QXp8vlJyWYCutMNYC01GwGPwBmVIqO0jZOLLpTocFa6PIgCMIJa
/IqWb+yFWKPKGwPjtclM3IRMEsnStvAFQ2Vh3AM+gMw8t8yQqx0i5MoEW21JDPbE
nU8BW2vsoJ9nukzooPTpbPP5UaIPaYBmdhAgo2Gm5G3mKsAYKFk1iA6LBxcfc25M
vBYFaFbi6UEBOKHOfnXpRKac4zuVSPlROgh37QRfNNH9/vRyi9t2JqGfo2fZDGnn
rVVF6Hpx2jB3o9QBiZ4am8ewAgTotlQcYSt+vdSd6Ec+mB4wYwAw6KqpuMYZvlgb
pq1v6IzRV1j+wbVR/U071rT89WeTfxZZ4KZ6EL7jhC6jxezhVyrP02tlisSTFNIA
0WetN1iY6lNHtprigXFq0Ji8Ff98gl7n9M5akXQonrZmcwyX2/OX8uc+i98sEilB
dqkBW9Yi4fegqNgP2lrfTprB3jp+ECtOy0RWWxC+7BCe+WbQsS1YapjrVIpUhY/Z
cwnqd7Pj0EjCodDu6lgOdIPYMPxI/3O4jYA8QVUSlPWtJwGvFP2Zyyku4YaF/8ox
yor47ypRUczoIgIxVaqfMIkYtD/KmpWZ79EXTtA9k/EAxMFml06goX0a/E/wQbLI
iYeFM62k5WVqrM/DQErWolRZ2sg2XVTSKDzioufMBYVGm0+xTMRnzhkOwXbm7vYw
kRuYiHGWot6OI1Le2CJR6+ZDEwlP+EcWIpnuVwqGg6PuU+c/N8zU89fQ8yW+w3DX
yYmHfopL+hQMSiC0xDvrZz+qdIyehrSv+UR0bZBChtr8urS1n70Py2Uph4NPni8O
HuSNiyM2G/c67YyaZqgyw9TX/psU0+EhwhtkwQIhd+UL/VhQkNS02lC2IwJ+/eq8
WVccpk9wYzP4Uu2s4VdLUllOC39B9hVhutn70Vta3CMv7scuygNfjMhZw1kOV9ll
2yBmA3Ghp5gbAx7ure2WC04twJ18zrgW/tpKtyE13VZkq0oImX0yOk1FfiKg+3gz
OD/+oC31dL4vHG2VbGV2z8R5kANihww53l4AloQ8c5CdZDE5SYtVgjc0p2rVm7P5
WmZhVnjjyfEyuaI+O/1ECAn+rB2Z1r0mhRFrwsvFBSX3mcYdO62c2uj4phkuhlaP
qDEzFV/EbVPQx3XcUKc9XP30SpebOFyxfC1QcO3WcKhCrtMrRtSUpm7aiZFYnX6y
4cIT9J/mPteTuP7dOf7X/lXwCXKLi+TRPi1dCkrWCt6L74FTvEF9FdR8kUlv8Y7W
VDWnHgqEH4cyYJLAdYBN5mGJ/bEPpTLLTZzjm7jKV+IcSF+G59ihfR2oDEJ3UYbM
J6OC4nWvpKuMeSbxOAeuKxSW6D7wfr2FLqu+rbXQJmzYm5a+vm6652eGpaahGt9C
9ue8QQx+nEfNbyuDqhwuVbdlvt9lHg096l1elDnsjdgmA7qKnOpHFYeWE/fMniXH
GAYZP/0cQGuJYgaqx3FW2LizB7ZngdL2s7L3A8LjUunQaE0cSeEmZV45o4JuIC+9
2/3NacvSIB2hIHxJfrigfIuWM8LF21X+Pd9UVbzR0da/8FTj0jThVdAhLvL3m4yn
rvo6Dla5lYhrNj+J0UJigkzbmpzrAQ3VRblWyjgALEmzXvVHbYWextYCjvV+66ss
sfwxMcXjmZLrkXhAtlZ4XFKMaXFYWjz2XyiRvbzSZCJKWK+pofd0xtg7lW0j/d6M
7Mo6MOoqWyltOY9BwmBF3BvvOXmnQe+bmQR2gTTxGnVzpuqF3I+PCUb3dlocCNjs
84O46gu9nCYTU52S5D8y+u+II/1Yp0VxiakQYttGPoDkLHfvjuNL1JTu1HSMvma3
O1fFkbVb4h6rhCgf4xoDv2blcN8WAhoG46k/VOw0X37/hFl/U8wfyIOAwtAyGn+K
e2U5aTlX2HVg/TCPA5JDyBc09Kd5zsX0B71ngBJsBNJphRTrDdE7ZKmcSEEAIWs/
guo7djsyaVV6YYO06sxt9XbbTjBw8e1fTxLDCM0KHPAhPI84xefWUlIzKwd4T3gu
Eu8dxiH7iXRdUXMdpCqdL3Oqa5E731ayOHa+KQs8fz/6O8MLVzL1yq1D/xmO0yKH
TgNakADkhwzsv+p1/yEsUm2VxN35fuzrPSv1lBBx/1IMT3xvJWXCsZv/9ODUDSdX
BS/j7yf5FQIw/zq7P+FpYeOMKK774JeBoUOvqZ3Zn/D1jcSQzmgobBMrQbanWJEu
utKqONkUAEzATs51Lemvhs5J5FBUCXK1kYw9jKyUtpgdfKgjKwXi1iACIugsVCCd
/S/KoMI2myq6OzWqLlVj64OQxAG46TzQQaXoicKMr6u60kzmGR0fA97R65INgoJm
eIOebrUhTgnuLSWyw1OCr2obaO0wyiDBAMFIQKN5gTtKNt5nd4E06+rmMHt91FGl
SVzyg7tHK+vyHCp5zrDYFpbIYzyS3gYDldI2XcVTCyhwdY4HnMwqxZb5wd6zHPGi
5TLUeCSEavMpCb+N573uKSBjCm6RHo7H82WCMSprhl0tDmjx37lYM1A4aUENyEJu
mWJ0jguMdxMAtuvRFXW6BFTcWhySsllDEtnmtYDOTh79XXZNdeOl3RoAp7JYONmt
QkeHhwTtMiUd7Puug7NEte3xId45GO5EUkxthqvRNda0f39s4R59P+Uobeb55pYq
2ONDziUJvJD2GAgwWUShUUHr19bYlXilfZHS9DwBvCP8i+rSCEiKNN58uc2w3ClD
P6d4rr+r5h8B4Ny9TGtkFNbMG+CiQ7yw+QXsh3SSVV4PotQ0xq1W0jKYuwqbnVZ5
++vduXQmSQD/2ddLC1icmBdyyGNhXhFTAslAJrCW/k9vZdA4Dr1GXq4EvuBinbDs
tMCaWMLIifbROUymQLRq5mmjOgL3VT39lQ/Fbm0Jvaq3JKMYQQ9NNcsP5n8IieOM
kwUOpRDcwmz8Wbc7rnlGrJExCDhuv+G1CyIJjFC6nwuwP0j2Zq1hmnY9AjWzvi3s
P5xU7bmcMDyN4YAUDdcNJZjxPj23F3YF0JiXVxxhJeFZgeUaF7lNPQNrrpkHLTwo
vJtw7qNQin5+wEslW+zQtaHnR5bUDXzw4Ad7s7snxi+W0rHddXbn+uBRyFfe5pSr
Ef3EVvKq4ei0VCsJL9oJ48Aj8Z0eApX81TUVFmuE9mqntvpc/jaU/DOzGdBOK/0P
8LeniHa6KuQWCiABJA8In0BR8KCZMX6UlxO7xQiRTcRd4Zl5z2onShHKIE5XqsKq
x/D0FP4ZMP04t1mghjKuM7VcnOiih4KJmFtTbG/ZU535ZEzrByhNAbytI5oY0qYf
RUAUseQL8O9TpUhbK56kySS12AXugGxbqEzrHOKQLw47ZwU4TLrlgRaAwm2iFE1o
4zwenJZ8apQ7vSTK5mq0vjwGRXTpDoZ04FhL7k+400aKo2WvexBLQMdvQkZCrDLG
pLjtwY8agCwJiuytEnjasow3e+0juRzLXYzMkzQFI98plnld0ygzhDHIdy6D6EZ9
FR1b6LMgEbbkEH//Om6vSXZ6Svpj3ySliNqX0DoS0mPDQU81SzXTSQie+tiWzm4x
uub+DffEs2xwv1+JVpA4qaLRXtZEvcig0C40gUWo0RrkpjwRmdM1ZULRKCqpuLCd
mjjBHSpNJv3fyE6z1Nh68/jtoIirKw5v9g1bQr4NBO74/Thi4mPcpMgv9n/5LFFJ
Ihsm1bCRu8EcyJSaaqCSZUGVIos5sQgOO+y26fUMLLsaewdjPJNxpqCnd3hLgV1V
8EV5LeyI28LkTisBtZk88t/+35nHylyXSFPNx3h3rxemNrxXvqHtUHp0UAzscP6R
gD/li0v6bEObGkIRg6xURyN+leggPBRdO7T+r7FH8m3YwY6QVk0vXjmVdebM1yTd
gtRmq5DQStHKvh9N/mz79X1GdRkNo8XqTt0hkj8uJn6OEOUCqImgj+seEV3NMCvJ
o58cNdGhbMYjJUwTZ0AzXiwxWIDV+XGCwQmzS9ssSwx5uIltzFr9PjrswZ51Hebg
EY+F8iAgC3lg4bpH6C2TXzpJ84dpcG9fgdLExhLRgwMB266mctNWw8A71Lfu32/i
U0scJL7D/XmFtjeyKn8uKrEyq+eSUsW1/E2X3ILnLWF9rmyh00D2Odpdlq18VycW
OxJuQ2OKHK/jt2wi7g+HkHHWR4uT+FGpxj6JUBx86p5Ug0TUpReI0NKMxwG9cfNC
gSSZCttQFhYiA5g5t6l59R6tdkGG26SN9etu2ijWg3/1PGQw3dDRHhQZ6zYocK9I
dPf90W+jVa8+GG21lZ91WTSh+JFJGHAVna0reRLXTfRWTgID0nbiesMCrVB8mimT
iFyBsVpr4aMGSnvSK5SxW/rXFcfHhvQkkeYfSgTeXEWzhh2wJ11KeOw9aoZMQ46H
rQLg8zn3I7SNQEcMQDlvfsqAPmLoWnijnJ0ZKynCKJp+BKPZgDAeeso7ROGcZfTe
i+Qxi/NL2Wj46b9Fh1iZ77oYfbmmb1azqnIkk+BlB4payKkBWfqExqVzxHE/ZLt5
JciZUAaHD93gmOozeFDXfUXDCYPVjueebyqwOGdFka0YXuY42QaOiPMTq6bXZ289
QYMCgZ/xrAnSx373q11qt6QfAyoEf8rAO6aBOC/Yjy0W6jE3hf8GoaR6hEm9R8v5
PxEE1SeyBU9h1vMB1JDw//qfZCUlJrYrlBlR8eWlpDBws3onGW1gEAiznUGS/mDj
D/hjs0/obxBsSQqQ9RujPw/fDcCKhrj8VTF4vWMoUnV5ttY+2v7iHdVh75zO3luD
fXysaWPR33lCvB0zFkbTXREUETWu5rJJSO/nXt58uAS5BlOEYv5HZ1jeE5qbZ0pr
4OACUyBmiNz4VyKlO7JAr/4QCRDoLuNQ2i9O+kPOqe9RxM3qFXp1fFohy3oJiYrF
cAcbpWlyrCd7Qylw1X9kXM5oDo4nymqTdHO9VWnGMZV0TE/fn8Q/f+1L5GUYKI4j
7y1Vrqb7YMd2XH8QoMCS7N2NjaNlZYXDj6SKj8fuQuA1bRJzL3uGB7PcwoivvIA5
6bst9DNvHIcw9IJGge3/bC2F0Pa5ai3FZh+s/UwDxJyvFOnhDQJiQC1TZ61uP03q
oyZCIEvo7VXzNLEJSKTzGuoIXUcVWYuvnXlrrLFgP7z5HLeuGvmmjcdslHKgzOpi
A3O/ak2HmN5OXA4sjchz8HILf0+K0KQvGbGy+O9j+3QF9lmSaivfnVaGJkzbnHFu
e4I5dF9kGfei190t8M7Nqz2Q0zop2EKfN+/P89LE0+G7uElc3Glqj4sWxBsvQgWC
uK461uMF1Po8YBtalMIsEIEtNq1exFwxcR4psnlR51YlEMO12ld2BjNaPhI+Nu9T
DSsYjBkvyHeWIfB+OALNu7WNVmDsY/cFBg3YNPnqh0uTq2L2FGv8HtPm+8IzMsJn
8pNCp3fuFyKhVUbGzo89ByLdZkqBzNLEXxvmdWCNwbn5m0jwzoRA2DtiaEJEiqVt
a4goSzJ1zvyVdM2l5xM5+hErcNc6SfF9V9Bn5B7JQz9QT2fA50yxZ0D15iRm6iHn
guNDJJ/394X0XT+b34ql960QfDp43eVHUqw9gFAjuXRrZMrU2puvYe5B8ydrE7Z3
RsY+L3jD1Gc7RkZYW7yEv+lLqOeqvoMrSTNmI7+atS/PcmMeS/4bURf5KnNsUzFA
ezytR/opsL1Uh5QnWC7lbeSIWzrGWzcqDRZHXiuq6G9jhN9mqwpjEkltia0bzV3m
FoXv/Zo/G76rzvkhEhzM5lS2xKjY1bJ5o1X5sHHWrDjf5xa3B8yoxZuw7XI+oj82
tc/z7mfNnQq6ZAkFCM+ZL21go0Er5c0wVvSkiiyWuwsy7QGWujwDzN1XhX/Qo+8T
jHigChmWIv6cpHhissB8FlkLWLW7ophEPLurB5/sn6NxGm3fW99TIHIiFodlJy4D
zGaaEf9cwVPlgCpXoeGUie8iUGVqpcoaPViXG/WP4Bbam8lHvBzHAeVqvZqkdMmw
N3CeTbsTrDM1VTyAl2joo3Bn9RclWUYYdQ5WXWDJJiw+XjpOnP/x+2XvEBlFKzSd
0gnWrMqYKJWXdCi/9bDjkNSmZVS2yZfmHz5upQJrw7RaF6m9nesGyReitcnnXI5o
SvzePMEE5bAj7CEkmU9SvVXt40n2BsnooUjdJRFDEK76ganEXst0iDjK6+VLZXUR
NVr5aKQ1U5EHVukjipjs2cpa0y0OE+S+Gr9ipVit2Y/W3jf8EbGIGNGuBaZT4wP2
lAAo06iCXnSqtQgxxeeshbJzJlVjp5TVXRbMYHlkkSmoa6wPkyEyrkUgIJe0QMg9
z4GWhsJI2PTj/A8WXY7g8oPZIT8qnwyym/sH+BgQ2reTwjyCcCenNrPqo0kKjun3
YXElGbafBKmwSJCcTu2rKGVh0AKKA/6CpNtEHWxqTnYiRTc0Vo59XIfXuekI+hJ3
IPM8IOt82NpzN854mz0fpLRRaWH4oYoknQpYEIreKH6i1B62YE5LtU9c/A3toTkz
TLhCunfw8cn9mudvfeYWLcYrSMHhJFuoCrOe9V+knBYuG+M5IUL3UVDzJhI4Lz8K
nwATcV7dA9aHlL/bZhPmPenyS315oAuzg46QoBUqVZKymNk0/FVj0SoQGAlUgGJm
HURcQHVLdmVl3QFqAQ3GK1J1cqeZbHVONJhH/MB4kkin4G4rHdGf2LkmG560fsJw
x4O0O5c4JorF/DFrsIDTBrhgfn4X3B8h2ZTnN33gX1+ML5Sb0FUG2O1lZJ3HKKiH
pqw+d/SVKbdViFmsIAN+DIrkKYdzNaJDlOVFFUsjFIq5F7QjuzylyFow3nvyywC2
1VUlCFjCd7LRMVEslDKKlTW1MD7MgUjwcelA+o7zrfGucvyCzvMOGA18ff7t2bv+
XDZwkBMvgZDCKAP47ZDdD+nrILQ3Y+lA9Xk9FJPI4lU3OYVlOPvk2UKypugklMGR
d63Viawpd6VK3wSS/kuQC1exKDIO06bNwaSSpQAsnMMkH3R3BWgkmnJYwaL9hbAD
ypzsSJZ5wEwyMeW8NJ4mOhFZv31+Y1TTAsYnzTG9x3i/Ibk/7Fr1Gep6K2jGEyTw
+vgEvO28WEClLAcOT5pY5mi3rG49kCtglfKGhdVvgdQ5+9QpSqF0hP2EBO89cXDL
Z6aZyHW13BU+X37LX6ur9dMlaG2KcujbBvv9mlt/N4G0D42Efb4a6PVd45QYMmfm
p3/0Ua+ZRojzXS7QAoY9Wku43pa65YSm1vV2ZDUqX44kIdDuBQAap7BslOBh9YtQ
f3y66DogssJkfLwIlGPsyMOh/O89332wYaE1Ilt89S70b+Naa8oxcoPyM9K2UbYR
FoKQC7By9B8jUcI2UjEVKhWqmYrezT8srtVBSYT80KQsi+W4bXy5uivZLKpjVIVV
jDXvc211pvOFXB+djYSCXNsgoo/gPlkfY1pzKbw3zEL5nCDRGxEqQtTcVZFe8HzI
N6w2DAwOa3TAYjjY2fUdi+o/89a7kdu1R4+23lndu8NRnBqbM7NcmyoSKBIZHmTK
+pZJKiQUMU+slkTfyMlP+M1zzdfTirGlGqwzCb2lHo+0idTB3oxY63TPKkv7F/le
3RTkc0AnElh8MmooJAtBZv2ioDPWz15GFhMmWoxbXM1gliW1HvsNDybb3e3xj+iC
4ulAEIRuktizyYJbTItpnSLPxM8TUk4WPmVZHpjpwW9tZIyIFBfb+IP+rUp5c1NZ
ff6zGiIz0tnOWsKvOoCxoVNIqyfo/lyPKFlxCaaZwUmWvL8XifMegYfXI+HSgpGO
8vgXNQTeeQCPq1cYB0YFdI+Brry8cUBcb5DMbEwNSxjwu75g/6AZcM+4nFNAuwht
15Bj64t9z7TLvCcjq74zo9vxKQ5sA0WMPgOEjam4Gzli+3Q+YYtpSQUAUPwJNgE/
3wrODQMkNBsumOnVFbPrvIyZctNbzH054RIn/NGvsBsLyST4XSAKexZ2569C32qH
IKi66ppGqnCldeF8eeFVOV/tYGjc5jdLQpDlPWtz/U/kUPhjDPRVr+f/o1XVD7lr
j65ggy4q42B93TQ7bNcVvbHJ/8S1V752S4MxVOCKuZIWDKebrV3uDBYq/c8MQikA
kvdfos+/Ku5wISwMUCUlX58GnOvG3jYXR7IH3D5SniEcTwgBwlc0tK/fSpkpTlJI
dJTXTf7PUjIzw9gnRZ4XXsdjOX/VTLjZxA8Aq5aVIrVxoG125Bxo9bZ5cmCBA6EF
sgceSvsLFnwNL5lVjm6dzytjDcC7nUz9+W6i3XdnpiuM838RTVnGl8tI2rml5kku
kW7Cx83Iu85771EbfHj6vg+9C+nXmUIslapAHFAAdidtll5vvzf1cKucWvC6YOs6
5DaxV4lsjTagCK79qNMryrhONO7y69G9cUiER1uMHvi5MREbESjBjNt8Fd+tI2dG
k/knzMPqsEi7km1563pZOw6i8vvGIxIeXuICE+rSe610zJMNVvqlFYaC8dXyFULJ
6YaRx8D7P9+fMfX5GDIrjvJ7Qw0SgYGed9pBHkLrVh7rcmyx4YjK4u858waPW5Jn
89j/8arQpkAFoJTbolIGgzIXDigollVRiNUbNIF3AriYYvHlhm3aTeUbq6ulAvRb
nuvUeO/zml/D36ZCpctEME2JAPyDF2LCWoysp0ZHKG8FN2xpHMRXQ69cIUEcSm+P
sJeAZGWCcKpK3tKU3EBhQyBNc0wz2Xnj4fykJD31IV2pllvp8tdjODWeWD77WPa6
P/c+Ft9Xma0dRepF3Ltfcz3SLheNsJ+UNYWkGvb1aQ2J1Ij+Zxm6GxSQdoe7N6Rl
BJHWHRHrjqJq5vlCvXvuITG51yvbnwcfdBUt7czovcQ/NVhjLc8hAwxiMV0QdIb0
MgVYOaMdjdDmiMDuCEDNj7xkTvkr0iKmVQN8+keZ3b8Jrt7j7LsDWHxW4s1X6dkV
wmVFdLKDrLCHkUgc3ko4m4z1jmiormphmOJKorh1XUm60HINsZuAqXJpdxrbw4ve
5yWHX+ox1QhCMPcU3uAUwlELBeNjzZmDNE/s7ZOaIGb6n3BA1SUDVrjskDM1TQbl
ZE1LzKnV4iCf4TGJKSsZdq1NIsH6GU07xspTAVnaNWMGi9r8aKhEf3vsmHnWPaJu
sp833Azm6SsuD74ll2k24Tw/uvIKK7Vrjth5Y4B3ZMML5kGqYS6VjfKtNGNyvbY9
syxExf25UpyNt+yoFo+t2qSGKDLXNqzXMRgvYgQAVKamNDFVRAumtmBoCho7qbVs
wRfqMTl84ZPyTEuwgLirw3Vbc+hl4rrYrD2ewmcw17ix5V+hFr6k6zSUo22PBMPo
JQrfFWLevY1ErMjikKxlDFoblqCbKfwo0LXHGWtVDy/D2CEVQo+kj8DZGfbp31Jr
mRKaFKwdQlI/v0/29v6ErSw7f5DGhcXyNeejWK31fY2e9pLZ4sNUMnEATLDzMYYz
FJFmDj5K9vacHFX53VCk6KMuLU2wX2V2v6+VpUPD8kMthfhMTSaRskgyjtSMEV9n
yPBTkc+jzrK2axkYI5tZyb2Hu5yH2TJ/Vl0BLEvY/04YAk5GTsuG8foCkjr7WYF1
0Cq3Brt7CBK5KHSszRJahN02WOsofOJKHAoK8Penb2hFvovi9ObqbKu5FQGwotWV
Q2A0VuVTT2uDFiRtho2ewsS0j6iC/oBNYpojsEkfpVCmCXJXMW4NOCspmLthPovh
ztn+hPfsCgomkzuHE4xHP8AUh0InzdUdVNwkd7l02gaIVv6dZDsS5NeGmUad9pXY
N3Sz/AehNdm0eLYEBMm1/Sy9f0rzp+/KXtcWnxaebhz/YvaRU0KEzJI755QRRGsV
HY+C4ESbh6a7AMw9760MB2fWRfOBaLfZzihPHWOdzw5XZEk7q29odd12aN6vPu84
ffweNzSu9NJtWRt0NJBChlgMyD5DK/oJjY5xFK4DZsZmijBFRvMcsMaW8z+mEO23
WaTCmaUN92lO8UIXZiEQumsprL5R9BRn6DFK8QbKl/JVTn0slHtfH8v8YBfyiEF2
B+eJ0zkaOs3WXzb8se7JYLIId9Z1UqnofFaSrQbqJQ3q2yjAgFtujdoSwc73S7if
HKNScN0pR9+F5sNFKKj5ybkilx7b0xHhXVHc5KSgIdApW4/gDEIgl9MUCXKmA1BQ
44Zq+rvkKXsoMHlWxFBSHASib4gNWNVQLIBbKGV1V1ugiLq4gEAZ/aq6G1dlwwUn
Whu8vHfNX9cMuF7Ugs+hzCat2HUa0vAlFK5Y3ROneykfqBdbsIbmRKxFR7nRV415
5nsu1cQTEMPUiO8PMyrgIdeiYcip43oGsgZy9XvFYkJuHNmCI6SotNxulhUecFdz
ExJGz8X43eQJW8LBBJyxrGiM9Q03//PKGwF+hkar2XMMSaL3LebUSYJPvmwXYXWf
FSLFz+tDWRzRGzCb4EWr7lDuXE2IQIC2kEcw0G2FObfLB+LsLxXBwOA+R1xEEEQu
s9BZwjsFAjiHUvAvgzu3M0t8FCKQmOUmAyJhRnAz4BlgzwlW1yS34HR5ja9tRVqO
fWIb37dVG5u7gavj0ZRypZduZhkrXemOnye4bze3R+dkhQy3Jfdw73rdOZHXtHMF
3q199MPkhF/RzIG8LoF5KskmANRbckLRCrpi6n2RnkspC87SC2cueWeLaIUDNk8o
FGIWusQUmA2Cc+djBWp3YduGNmaV844bda+Vsm02G/Eni1/DBJGAXLPRhZoco52p
Aaiugq3W7JDmOe92vC8d5UJIdyKaZxUEA0u6XuEdr1eGC7G0StxUVFvlQt/Mf/lh
vqsq46iwEpT2RqY6DQaboLDMcWKguvWS7AVNUSwqcyHdN1f/IkBF/aHkqIhnWoy+
vxylQT54f25tJ34aiFC5bVxngB6oSHfMZbhB7Hon7/EE4HD9Qo5L9/3Mqck/cFxF
ScVnU1rxegzfSW7TtOtOnxznNdzKmuIfwGMGtJXRdj1G0jIhSo1PvO6fq25DUbS0
jkDt50z+fRVxtg8RN6xBB6Oh3RaBNieOVo1vQSSuZn6e4YBx05rMyzSs7d9TCIAJ
lQj5+k6ZhERcgyPlUJvzSfrZIGEOAR7E+ducg0VuYDQ4ubrxQiDzVbSee1n7X2fu
OGPRCMmDLTROiW8nnQ4C10ay3vTBFtSi+9hfd75PM+AOOqiCW5FJh71Dzsv7P1W5
azYFaNCANbRRRR4raCtmlx4HyRqwb/Wt2kGAih8Pcov4o3PqE23yMXBojokofvgs
1kqteAdE/ta7cLyF91Wn7zSShr8Pijx/Ovzx56W7w/6uDypgsOdoY59evF6+bVbG
P5uTcSUEABSxqvycC1kO2JUlnwx8SRboOEE5J066U7bncXsEsTI7leBw5Ig92Pwg
I3+frfveSs/Z/zVpyiI+SIxrWlALzmljOzSXqHVMLRe8N2NCjIite857r8n7BIKu
E/+qsWxxwkZnLh14kFnCBBNooixY+UUofRM6grV4gXvQWVXRjnPDkqsjx6jYwphh
2O3HaZOp6L3Kz+GeOtY8D80pnrcLi+GIvzqy+fRyI5v9VvXEfm7aaM3TO4tgRU+2
RU0EjUQNrGxCog6T1nMvwETJpR5tyJsf92RV/QnlnbuKYIPyK5CFgo+TR7hKdaPh
LY403QNM67GocOHTNLVJsZBI9ih/MpzYQYqDXjQv2GpadFozki3f/RGJo4OtKVLT
I3d2XvxcNi10x+wiarltb9RntSQ0Za3Bbg2l+dRv0Nm6RSkkOcHXnzN03wpgPcfh
T4Lva0B9lvD1C6+gFvKl543u5YmG/FTZuyV7DKOLIO+ZFZ1dn/00tWezTW2JLbzX
amPIOrFFEqUUOajI/pEfTU0K5Fd/LZj8pw8XU0KI1YtpZe3qqY3CamtRKDpqBex/
ZBhsrMLR8yAMiEoYLP0VvL5h2p97D4scscfgJWDjTRIP3tC7tqn9NQY+t2mWPd8y
dH/pnJTUHm2xWfBbFZjRIdxwWSi0gmPtBdq43LyIP6WIHpcqAGxEFAvx5KkkoVna
AR6u+T6MgWcLpB8H9QQhc1+psNQKOIt1r0kJJIl7QXXMQpsovP7fMmW2iYY+Kinr
MJKNlqygamJjtMofdXTaTk3Je/9Yopl3nV1yl0uarkDN5bnEjMfyaJCDWreFywMi
FXzfjL5fT8qc8mBtr1YGs2otNU7eHywvTkd4Eek33kut59HyLeyjpv9anAlTaw2V
MOArPAva8SJQq2jlRXSbaGcpbWHXMUyi8I4gq8c4XlWpdBJ3A44bMoTjyIySRGwg
Q7OWq+CnAaiERV2GboLYsUwBN53BMPy51c4mGMPCJApxE3tUF8ZTwpj8Wgnz5AnX
kpGYvWu1DXTnTmUeGokIHy4f4OJPeoB/yJeBX2QepzKnE5FTvYgzbG6Z8GuUV+c6
ceMH+wdtyeLYot9YVxiZ+Y4rvnU0Fja/TR95cBnr1dlhKeSCOEQOrl5zO+yZjves
EwsvGCyFjILXiH6GrY4qwRnx8mjXF3mDouAkfxXla7072c0ykpy/hF81qWm8tAmL
NEr6YaiB1Ntcy9YaVdpi17Ls4TPLyKOsqe4HQKV9ek1xqllMJGQStskeQSgJu2dC
TnpDol0+xCoh+ENt8KH/bBYi8KHqOoKV6LkFYogmpLqPvZ8cZPvxr+/WcpP0wWVH
N7MzHjDcnAZxS+4UmayaOHukWlMLbkfs1Q4C6S9lJ4S+AlyfH/66HscIIIBn4lyY
vJbTJAgDFFk3jNv916XVzPs5rwUxql1K+FmC1vo3jeDjZ+kDRhjBEaVHDOIC314e
oKpeEOXWemrZbiivO+m5T9FlESqomPT2biRMr6D+JSf+vqfNQ82A7vUkYcguiJvA
WYXyE1jooqsrPMey9BK0zI4tBnmTkPKOZwtqR1Yz0OhBagAz+7IFV7FoBAziTwCg
wQCh+QKLSWug3s34g63x68YCnL8iK7ilWyAhzY7d2WoLVIySBYg3GAnSJ6vJvvCc
cLX9w51pODOB6/T31FjsKiqSdhGvCoRaTzSeJOqk2T8RgAbc1HDH4Rl8esB6fsAQ
oS+eqpcO7cRZekhWRm7QAJedGZp8zl5ByYCLsfZbdww50yl+eqegYQBv8uxqh/9o
km4MhsTQNrFFD/cwOX+cvn2WCOcOnXM6DNhRG3sPKCbDwpDWqta+xDVoQpY0XBVJ
JHwvvm5n7b0QDLS+zkiYE5iUwOSut6h3f1goyBhkmtbdAWPqxiCb/wj6BG41PT8u
KZf6210jGVgwotoeqRjcs45k5i2Tx2mAwXfBxXkRMfL6CThla359SFciijTz4JMT
wTWIVl18DB6/i0XM91KjkyIQVnPoIL/Bz817qTadRNV4QCSmw+yrnOnS0uPgvHRg
6CarB+qr7P4LPLZqcZFsfJElzFIvtvKUjkNvnm1k9gKROT4Xweg9XuDzfDxGPpt+
b/vWBBW0TSpPjmIaTQShfP84ZmfyF8HiSFSAHiALfLWmzCznrJDJ9is4ONZf20E0
nDzKeSwAW84fgWW6Bq9NsYYwtcJdFPhY2eRAFSIstLDSDaNupid4JVZ2BMD/0rDz
Ia5f99imz9O4UbT6p6Hj+TNsGwwXZsVweBexrQJgWigE2/eoBp/xSj5wEZqFyI1o
2U5JlMgtmuiLrej8+EDMPfKxOeZjLyM4/K2IpKK9AJOuTR//o/qTHitP+6Qm4Xpq
gCDl7stGSYxgvTVmIU9jnHFCkDUJlCmsdL0R0BgWzJsW3ILUr8ufztdmfvnlHksA
w8c7eVs0s4ZEJkb9sDteKvkv1cIfx9Sooa/0gksnzHVFfCd9cFzKBik8GcZEcRGA
KVBTsxdHqb33fEhOZMok5r9Z7u6+8WfNP1jMxOrwE0gMvmvjhC1wQDc2lqInJVYu
fQHLmI8lkeye/mSwXqOgc33bXoZLWheSc1p+3LDwitK4oS+oUm7OeWPQR0MwvDY9
t9GW3C8G3aVN9CUCngra3CEKNf4aCFiyeN12FF1G0Z4vMgRZIB2fQk0OW5Q/8qmr
PIEXuKLeyJaNi+73/Y53pX5tprEBryuCA5srUr83zkCPa3VsOEBQp0A3OgvX1u1S
RE3kNdYAZEoJh9avrdPdT36o3HWh+iFW4999Or1hu96TYo6GfDgMnFKnGnVl6m0k
66vksiFCT1RarxHCQF13MFHIcW7Gg4Yj2YoRKoNUJSY6L6trLuMxxuAxk7hA14DC

//pragma protect end_data_block
//pragma protect digest_block
R7sidc0WzYXviW1WUhKIx9TQSIA=
//pragma protect end_digest_block
//pragma protect end_protected
