//__ACDS_USER_COMMENT__ (C) 2001-2023 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
//__ACDS_USER_COMMENT__ ACDS 22.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
j/bD0x/hewlYJ7rQuEa4K9+uRJLSQgXTuWLSDT4FTl46bZc3HJKnGtn9wlnUHWmh
7KvymwO+QrJ8KhvupL21sPAovh+b2tJj+PbPDbXlwTw5Ca0L/j8waujjZUmf8wr1
dtGpI0iD0aeV8Cc5lgdxo2JHnrPMsoAvJQ/bWjoiqN0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 11488 )
`pragma protect data_block
rqBH07qDAsfM2nNsfr++/LcoN1zHwMFCv89fx8oAnAPHNU8jhQM+kTAWJuI89+FL
uZiQkfjQDlxGKkYszljjCmUMl2y1QlfAW2Y5tuu1OXMN5LjgJkQBHHSIxr7mymxG
RsIMlTCQaIXUve54W7LB9ZvLPw0jxRAcLcBrBxzEZQhlPru4zihpK38KJRpwXQdS
eRsc3M7+/9ioTHPoXNePF0qQCFlIi+Z3vJgrD08ta5TzBYQxm6WmG5QPH0Hyx0LG
Fo2aMbqEqMLHt979uvP6lNJZ2Ff0PqGZa0xS4JyGusaOqODrJxN7IU0WitZZs8M0
54b90Xy+xfQ5Y0lBEkaAl/km7g5Bli44oqopGKzbzNU+Lk0Ru1mgKT4jkDGLIAzp
nEjmBf4xH6HxS4HFBpe5StlxMdNWNmfFOIp/jd2wFnn35B22R/o1kJZf02cmdaKu
cjCFCzmF3vK1hLK8aAIMaL2WM5twHHpZya6yJCguQyaXqJ0jsC1gfWxWm2nKm5bm
uPHNP8U7pkQ3URXFcaHmCGWlNVd9xWzH3EUh7zpmu2GhnOQyrPUw8X2IPF8XSXPp
4M5lcgRrBp8UKAcuiKiI4QfAQuyYozEKjYSoUeJXNuCrsKuKEBZuTvPyc3xw2Hu0
WEGpkXxBAtG2lJ9J5c4z0T3B1eCRW+th0Z2JNe+P49NpPXLY5lJMUHbFtgh/i0Tl
tngHUvvFz11Dn6noYtAZA9mOdrc3bzotkTYXIX6qLKzbvEeOt8M2zfamh6pKHCC4
rKLnTp+nBL/Fq+lSi4iAgrhb0Q2K5NVNDUp2psZGVwzPFPDXqAIMJxIKZqCWiMTX
08PXTccvaKhl3aZ122QNFLCSqpOqQT3uWdB7u1Rk60cwitvPvnue/815+ghr4ztV
srwgqj9fGrB8iHS9KTUvEBREPuB/QigPK9QIqtEOPXSrPPkSuhXYlfLQTYa2o6BI
PgCApAdfFRUtJEp8dYuSNe2oLqljbHJwL3cTlsuzdMkrFq44pLWYyhCx6Tlm2C2r
4I3J5GZ9wvoXEVe6UsFoKrP3nF5tv/pMxj6WdGvVFrqDUgWtxj16AN6AAM0M47sC
5LhOEIMCYkXu7M53VCNdEfS1pRk82FKFaVdZQhgJnKBiVHjiDEmfKrcQCP6eCwSd
xcabqhj45TOvMbuRoYk2hWvku4XQoEQlqAtBL/cP2Q89ihBVfB+i0PgSY6V1TaPt
/BFHL6pxedJMVK02sDe6wVTjFhNO2gNQxy8xLCQSSIFo9uyC9ZD4tLvNUkl/Sxim
S5JHVDaG+dImLopKxK0Wdo/4XVSXjbW4IbWl02Er7W9dl381cZeydvOev+Lw9n3i
19g5uk0snDpjzF/VI21+wB16WtkgxigTKnqXUp+ru+MBeZnOMzJv5/vMs8MwFsDS
oCaqYA26juvv2Sv1kx78i+lWi0bymnr34VBD0kSPg0QRtmS2qnOj1DsZ+w4HMO7I
NU2phfkMVpMnt+/6R4fotSPVH/fw56pEhaQakabMQhLf1wi1K8TqIVReXSmOeeRv
A5PR3JFyicyKP7w94tcy16ffBqHkuPkD6FJjz+wA9UmRckOnDfElXfwdAhybDGgU
GQhU0cljJsUEmjlMroMiD9p4gnZc1iDBMx8LI0hE+n+1G5QkAIi40ZJRqAEdEw+0
QD6mZlwtZFRNQwTXFhTri6rtW55DREXB4Ue9UFZa6zS/ZKqazAXkMmJCrWGfqiTs
eDi692htXgHYDruAn4sbvL9itnsTlyN3oEDTpFrjBo5zVXCn2SQhJtyGNO/2Q2BR
CLG2Y5dTHepiRLUtyqdFCgq1uW9aw//Sstq7nF6QFiTlJTjfrYl5UNNJTSxXyqT3
VnB4fsesmhgC16NJQIT1q5s4MWZ7mBXJc6/96ZeiCp2jC4VaxgsoG2R+230EKNd6
KruVw4WGoYLeWNvYKfIm/DE4tXYcGIGUar++gVqr3IGue72taQi84RhvrrxkkW2A
+ItA2OUfQW0CprC8nGy7baLnA3S/jUx2xRbJiPafbeSdfLU89i0mH8thxlRnta+v
wYtiT55zxqIa7Plr/TmWijh178KvHOZpRQmozItjfgj+LYsRFD4SI0eROJbZS9fx
cAAOUlYXSXpJs9KgY6i58EZBURHhfLzjRbwWLUrMqC4WYZAnPrdAkf17rscWsVea
qdogWl8bVVZbnd80LvpQrS40ojG2ZM+Uum6Zdghtzd2sAEZU7h6z/Cy9XpBZmwpC
UnoWNxi9AROf2IhQfb/KSsBHX+KMsxepxSbAKWw/Rx2zuF1RbDgQ94jz8L8eydq4
USpaJOkrrrdjkO7NMYIbfoAPiDGySKbWXYS3WPIQP4w74aR6WBEsa03Y/umYMA7Q
tC3SXtjFm4RkDjFK1P31E0dNtnOrXEZhXhwoFMigAu9MSc414QDRJWtK08kKDKsn
g8ttJqGQi0LPJyQlnzE9A1T+0NtdEmMogOXUzqw8zMWOj0pe+l68e2gFH+Jq1mzT
Fty8W2BzhFQvA0crsfvquDF97LgT2JBKeUQT4FNSGW/cqAhmrFY2vKSmj+LP3/5K
uRFkOM1Oe6NOgbpmIXlx/Lr5KVJzZjK4wWSf7x5rMyXKWCJTm4IzWTyxW9o4WQ1K
xbvpjWqHl7OBPlNcJHhxVZoOQFPNplk9zjYOKMNQxSbAgQJo3lGj2Omr6q1/VwNY
kjRijzLQExVHVL8pLwUyVoaR0w0En+jRt8yxNo3Wn/N5JXySBLFieWUgacnVf97S
Z4BwNo0/yPpxyCNNGLC9cU4MCXGM/hw7PLcIhh5fTvmr1ebbAELWlW6fnRhf00tM
6PGMaYdjvOvcrHO1i8iM5HX/PxuD4Xc/RJE1MMNaEx3crxRyRgefL4+gPmsuzRZD
kWy1JretIUozpU3u6PLupBcD7diVi9uW1pTWClYW28aLLrN5i50wdJYS0l22RRQk
rwPQATddB9ujp4KpI8ycML7A9xs/cCNgmbBOHDWQb1h+q7ou0HwjHtk7Y//a8WTh
6KgCrp+t0JpZnitA6wh/zMaU+K/ndmWVxIYDfV1RaMAKaHwVJWwDlgCZv0UpN1qs
yFDLR3pj72X0htwGvCIrPbDmGhnamq93CafI0tik0zeTLYTFpC3rRBBmyatC6OBU
hJPibvJfSR/TZPINg+NzjS4KxHjtf1v+tmCUXJHcROmk+cAC3dU1yJPZvSsGS/yC
eCaKTdEFho8JLebKqz1+TyM7D0Xe+MyJmokrgzedSCPbviahPHqzHHB/dAGaj4iU
Eh7QLnxsiO5V5qsUpaVFxkkb15JYRDIm8S8DU0wQ0u5BXa4Y3eHzI6ChQyvWqjsC
0x5rExnkMl62dKuPESol348ZEKfYKhI5olGyWTu9TTugFCnmf9a0ZxCSp5j4Ibq0
AqjuzaZsZo9HuzY2O6QoTYvSitkcuxs2AhMlyhGCYASxb7eQA/h032uJfjh/27zl
6KflDtq42w6AHCz1clTzNUGaYUnJMOPpflDzHFi8+SuRl/bzx7AruEAAR1f1l2os
uqVVhXhkBaJDEssD+qxedSodYqouTLBgWHuOyTlmeNfZl+Uma3lPjXUtz5ONwd6m
X3aeWPShZCcXdsO4G+FC0bH+PbrHmRoqVSxn+w8zr5edbSmkIoLiVWk+AptAClq6
MEykBLhLrZs/t5dImN8g9UMzp4biWgVJZoGsrX9PhStGZiYJ6IXZ7dcgGS+/em6P
q1phM+DEkWYcWqcM6yf50vKNahWD0ynhafNFxHB3nuVjYcAsW6iMcf9AGIjCEM2A
iIAhdAYpI36ahTk3PdUqlg63CBCt3OIlOrN7LBJJGY7Lsq5ZzDdfQL/H89gGOd7e
yQ2u7RtmYPnj411NUDihiKL8mPOK/j5EZGFb+eU/EwDhB59FCM3Qm3pMcxQZPg1R
1g2G7UgAY9OR8tTuP9PzkIBybimJ5MA6I+WeepSUsk06pEEQzbeDThCIlhfz6IfB
6gsCJQtN136/vaXVJR2SRMWzCMlsRECmANfy8h6egnk0s4DL1OCcIsh+fyiWVAuS
SvG8JLnz2wh+YAj7OmhpWBgg2SoxY++JgX6dWRXvLs285nBZktyocOg3HNqOIumz
8u1eOP61rkm2ZxRc+OGKvBsVvAOPgUTTClFLkOj5UhqNGSvj91nABM4NkgKgARU/
HGZJbWDiwrxhZbVrfs6q+g8Uyii7LlfiE01ElVBLIPx6Y3NiGHR4BqRfOJKuqVNd
HBob/T6220X9OPraBMQH+o7htJTqDKSjr6VMXlta0pRxJXbq8qoDdL0cmEdHzoGm
X2Kzmrlk2zQONqViL9UgKJ0dOyKLmIxA5rFgCIcRn8o+m6T+VZfO0An4RrW9nToO
wXj7ghEbM3pDpPp1PWMLo6sSJtzshjfl6rVXSc5rglWLN7c361D0zEX1zSzDQc04
PhOMWg1yAR748o3yB6eQs8psaKuaFP/ZNd9TWVMvkZLk0NyIunDby8+/HBuyXQAR
ptkt7Z6v1VPGFe+rGOTZ4oxoZDRcNgS1OiBowfPXdvGnEdLBIz0BZvtbVdDK2biA
/Ic/ZZumwfZNpOYnbw83PbU/Caq2YR/algrKeDopQ5fvNdnJldKrp4zaTGxD0WRG
Ah/TUfN+JGqfBKZ2UvtCkMj92fEoHbETOR3vrqLaQq5GaKRyjnIDZqNs34B0AEUj
kv/+anvyCm3QuJbRh5H4I064Y33di5qUlO6X0fztYhdqe4V50aJgMkVAoA22pgik
0V4/XQdvvv4uEITgq/aPYTxQQNEpB24ZV4o5mvbrkWsAn9oO6rjCjpBxJ0INuKxt
FOzOX/nCQ4HwNBrpIh269FUKrvThqov6zPTM2Sx2yoYm/pCOtUtnvGvnJtsoJ1FA
maLefPgnfLHgOkMjpaYyzoKbgIEpa669wLOFJp3g5Za7kG1Q2ycO2+yl/Pfuk890
rAqA6FSBKOyOy/AfxjDRFdsvBkSlpbLUEVmyerBj7NFWSPZmPgTNxKu965L0njhB
/mbBTbF73G9dENO+bXXjLHXKZBsxDYpPgH38Ihr9OBw8QMldleJsA+YCDo3wyInw
z72l2L21ZyglBJP4Nx7/bZTNWOIp39Fggi4i8DXdM12cZob/F3wPn+2+VFbB6l1S
QNmyVG+YDvIsndhb+FWdEx4+IKcb75kRIX38ppGr8xrPyKEgsZk26AtagOaspPE6
HK/9pjBobxXEnn8ccPLffq4tt2bkgvJvRswUDgP18Ath180g2Y1XjpEEkXbsnAEC
29wbmIhOFk9zgXaA/Sij9WzTxQFCUFtwVLIjgS3IU90Q9q7TvkRiqBTZR8cQ6klm
UdBKuTG6MBuGpS4LsRoAYC8Shg0aR2x9K907TQPrY8dw+1ySKkmhADHpHqB82d5N
BhsQXDR6871jb83NXzksNQp/ECIU+emKzdp+QkZGrglL53NjEhDz5UiHST4qHoip
aOdFp1q9mH0p5aLxy7vga8J9Q77jJ5DxBrv0iTwO63bMA6mw4rfxoz8NcUoJhTC8
xvFQfvSIJqVmJ3+9SsGvCxlIBdiOyDyPfoeZmJV936ckg1JHEqoq4ubaNPEBtAOj
0dDxZ+UXomLnQQicUDwQ5ZWUx5xqeryNQWA5WZKcqFBftvbdTX5Myxz/PbkUya41
dAS7o4hMvfiF3+TiaY3uDHanMOdXwFAnZbZWTOX/5C/iFs+luZKtYbqY3n3u9683
kQDJ/Ms1x9XmzXgDzw+uh0FXpvbNUhfesvtqYjsL16EbYRgYnjE+MsEJ8/FDaALU
3mEnFzTDxceyGZWEhYgd3N9DEROmfnDgqFqcoaihMwri6XsOZnEwMN94SWyM8WHh
1fhpkk0Vc9/GS7dAImBI2LM8+DcPwpVXJ3RJJucUOZ1p+IXFIgDVnQK7M3ybcd4l
hCQo52XIdd8dMmqxLbWc++tWLARN6+gjzSYLVTUlPsobGl31sGAyTBbnase90nN8
mXkdXg50M2scq4iuMeY+NK7WvmrllTebWi4lee169HrftC2XjQFntXhzRpUtGnqF
RdTWjky21OqcAWpVV7XxBDb1YqzS05kAJD2wI2qkvEs5glGP2bkvNO3vgKyAhQjL
KLU2cc+QjyATVYJ7PaTQQyCBJywdaCC0ZtOQW9ltzRCV4cT7Tw/YySHGrzBmwwzR
od0JbBvwdtHb5jdrxehJRo8LjxNibs9hLftoTC48h8QiNtKZW1Z70as7Ubb5NeSQ
tu3/JR5vpboKQB85CCHS+u38tZlgGkyYT5Z1u7dQbpAl6iUyJ1V7Fmkbhg64GEUn
e9cu0F7GlcC/NtUu20p6xl9pokQxJncjstgDvygY5MmFw9ohVuN1OzUeLbMzqCyk
wSPnTftHBAUtdqz+HUMP1M/TfF0MAAl1nj7XuY1z/dL5nv0HgVwM/OJiHfE33wQM
gON2SRCKZPB8oz4Q+rPCNtdPaFVbrQqjCbrKaVXKn2d9ciaDA6zvTJK8PxmDr7hP
nOsDRB9xDtku9zHy2Iq4QBSaqC1wk9jH6tXqgNIXb3CbF1aPUhSeBppIZiePP/i5
LCXdmVPekmc21bcqZMqnRO22EcWLafY6wuU0ZtmGGSsnVirLbrtcw+A7geUe8O+Q
sP0fJog9f2ehmrUhlClTLRn3OVsJSEnE66p0pQKk+tDeivBtM0m9vL27GfdZ++Zh
9sML2J460eZq6KqwaoGr01VkUHij6JMkcoIFJtEkt6jvPVVaN+diBWrKjA0S3XN5
qwTqorgWnzO6cjduTi9jbLR1bErOfeZNVzhSI+Th+zUUf0oL9lZ4zfRVQmonYiPK
3mYDR2ffplanYFuVwZZB+grxlU+LA+Y8eFw+Uo7RHj7i+xR1koAZi5kEVUQwKLJg
pV4w042AjQ/Cy8OyZjS6BaCbqacuYmElGGkWpjbNNJS9P4CPRnh8gILFhfwEY2Mi
y/Z+Ds6MwcRnFTIm6usSS4DvinsGhwxXOTvza5F7P/R65g4Qy8tJV+m2u+247fbh
RDijVUstzGxuzVq1p3vJmlg5dOcJ/NsfSWZKQjTtcDWNMuw5WatLpMy95/1LK5NF
ZmGAMEwbalhqy/4eMy9SSZmn9p/V5KYz9WTAczKliNQXptdZr/0xHP5H+s1mR14u
6OKJjgO2mWKMPfvZ8bbVObM0NMS4mkRLMvsUecVyi8iG9qpz+qUfXJhMNHiTsQZf
HigEIAVnuaoIT7Xfm8ZrdGiv47ptTPVsEXmS8VmybTtOgzRbv0cC9kfNnTNw2/WT
4jpNr7uILsN/VjndecoasLrCg15BW7fqiJvYeOl6pViE0t/iYn0Zi/72VXMyzjII
wRX4WN8cqMk3zbom+gaJpnnLVrdc+cWfiMPw1RQ5Av878L3kdsIrhg+qDCR0Ur8L
LcDv30KCc9rHlzh/D5got5mtibBbcg7QLdPbi1Z8dClaz2Z6lk8RHiL4Yu7v2jSk
LrTasfJSMrkWCUwnw445jip1V8LpJIvWBLCxiqXq0nKDS3Wj9/qguFItRQw/Etch
i9K2AyE4PrG2GM5pFLyCY88pizZ3XcUroNyZYFT0Usv6RknzU0f2ugvRLG1YyqxX
2nGEWHzvUm9E8bMOipaBg0WJT1V72EIJwWPmyXJxcAK5HTTBfogbLLdGj/qUGct8
CBaumRnwYkSLMDB09r740iTYyoacgrX+HKQ28xD9w+SBPjsh4GCVO3j/aNEXRjwv
cUUVbGo9xgXIa/QtOo0C4ct2FXZ+fuqzu7UId7bLqzvKGPAoyq4x1JYqRCu0uWiv
MlpVEqfJX4ei2XrXP/C6yw5hPvQIcoIG8GvsZaVRdO9X6e2i/Qidb+PvtDrFS0kx
8pnPNdj9HkmimMWDjIoIhMwo7UQOm48RWBUle2mhjPNjefxLuBwIoJhd9QRT1Yjw
5wEDAwhIH5f1UJmLMrqc032Twl13Xy6prrWERKEwyEzkhzUf5AVRdlj0W0B/+eaF
9/v87k/s5SOQdaCwR8awZ2coeINbGchfsmRAS6g5479hBNbBz3CkxCeJIwjScn2C
DijIne28xdLwBCjs0vxiFwhn2d7xQteljR3uNRYtCbrRJulzzBAYk38KCzEb1Zms
lcEiaN6Q+BRwotFneJmVJLVoPuhcVuUIEYnQyaFM7IMUxMn+ZPQAknJiZt5drU1b
TGW0OP7Ovd2m2fQ/9vbScKgbteJKfM7SvI3XaJpb5mpAHIet1bWh+eJyUTxL7HUJ
kfMlgY9w6WjKrW9nd2MWzlkAyyCyIRa2mdUcu9Rr9ue2Fivp+VBhal8SYLQeobUH
sp4++BE8Z1+db6MPFLJm81jHcr62omXOsVTTezGUP5wwH128whu+6j+fh1zACyEU
NTCiikGwUtc3ytaVXU0pUVFjA1uqgqNztSAwCc0AiRW3ZpgwCgEefiwgQikVYSfr
bXTWNWyXr4Nf7owIlnLoAKQr2TCDM4vFbwD4LPd8IslFDblsccBZdIr1rIKrs0hT
6ASVVx4X1BIdQhe/gA3u0/PbX13tX+uz0EYz7ICs2JesEWzPpbaIshWTeWB6bdPP
tjw+8k++l56P9pk6AEIXk7taeiuHfnYdEm3oaG4QgHU/AeLXiIPFz5N9Smeibkdn
yDAaj8GSTYaAnXzUO47mslezr46zN+n6lX1J3G4TtiZjghhE9aMSxgCilCMvLCuE
gR5O/HYCGtGAn/PLugLSTdzsEJYAa18ky1Preb3swUz+H21drjO4cML6G2sjr83g
gQmEJ2LJEfmSy1a8XCezy7R5Ceh1ihezTQDIipEYKR/q9NAw8aRiKxnIaCgZ081m
QoAru0TZuvoZA/M5wDeTD618URwezWTPItZbaqX7rTsipEDMnq91slGrBIpwH5Kl
oILkv/HbKL0JScPRmdDCZ127vQpc/hhNmmixtl58v2WAJXFu1cCvEcqOTORFkVhO
YZ9gkInSRHX2sC1W+92eq7mazmA4/XsUaJIL1ZS0crhRxD6QlToQaOE/7FPoq6bN
r/xNteW8i4hXxBBiHhxOhzN1ItBWZxLL+KZ/EWUtGPEe9KrV+JmImNip7YyrNCuS
GTiSDhxhhAN+JVjlncLm5gzzgpIkwPSEO4o2ITLffoSnRLu2xeJWOTwbjG830wym
sHJRP6slbyGgCxIDapZFIHu2vKw7TyZuXGuJTGW3JNWCEb7SRfpPsUVqC/+Ylubc
kc3mfhF3W+5Vj9srr2TAx8c+5QuxNvF12mR8CJx8lMLTWFe0zRDdRHaVSRRZ6/fH
jAdRnSH4DRqB83GZ55bfyGn/T7+lis9wjtMXaX/7K6jn6yETEbItC47lUYRR1YGU
+0EIDiZik5lX3qV1YG0KU6Rf4gsxgVMCTQbsbqEh6tM9cqK385ybG07SbpXEUiIT
QUZvN/tMLGFoN8nQq4Q6PKAKy6OzdaP1NL/Na0MDqNGYNUdyfRj2ygD1t0UqOfAB
yGyqMWoXWI8HFSoOhMPrNEKHz7GWSsdMW6iY/YgoKJGumZLHrcLVd3CE4wPqee+5
B4wDRlSD2we+3oQOeIg4JGhxU6xFHlatJvGUUQwge7bOrLVEeOo0APdiyPDOW1m+
/6tPBWHEo1PAbUQkwY+qNoyUaNGoFIYGYNle1JRuPjb3d6TuFcHF1nLoBhmnCsWV
iZbuta2GnjWdSGC5Zp6trer/dP0S+nDkYFMnwvjKu2t/2N43TR+SlDbtRQeud3W+
ONLWiDPl6cSenRYGJwbpycuaTyQJMaOsGOisx9vgSsnSk9fxvq3/3FwEoJeU5ABR
NheYgaixfmPCR96eDNvmDKWXhem+FHioP2RCdK5IoMBovYkwMnF04Jv4cRpVn1Dc
iys7Zp364qlgu0LxgnhwGSI+/HgTjavkLji+nNt4uXU4+WWkjFV7af2aiAM09fj3
zTsNk97J/WRrgpgZNCjbWTtx+wp/EOaUkNvPt5A23bUwoD7yDov6m7Rn/KNV6gLU
NqFOBgDjqLc+IO6BoPx7Zi7my516y9KHZXK/E/2Ph3XeyC3rBRFUi9hEJ6NMKLZO
q86MTOZsii3TlQ8xSDD+f2GS8MW6Wckx0zWF3SI6iJd/l338K31WwJ9aLnWdeIeq
rdwgLjkdITcgXtfy/q0V9kRNr60I/VFUOChIRCm+UNEpXa421T011qt0ZRt/x1MX
HQdVlFI3NLOxYomV9bVQQKDG4AUocKZU6Dzu7i2XleIQ8KScCd5CB2TMFm2X8Vgy
M/aF2cgbRnwL3Enw8mySsN+wEumCe69T2FQovEyeZcWWVRCzR7i2hqDWJjxShyBQ
SGJxaNindszWowUJtUCjn5XUFdkqVXG4octiQFs1i7pC3KRI4Qn466FMp1r27FnO
pkO4Cz0W1c9oaIgE3OQ9Fq323XRMZg4EbyKW8OiPqMv3cvXmujgyGM8CgF9lqtIm
VtO5Gw7sZpWOn+MgCPIm8VNNC284r86lqDcx1OXBFAUcWX32RFLWMm60JsMsH11r
LP6EBOI7ntRk7XvqaR/hctOv04W/a2AHj0KXKV2YU++WpKmhRFNyEdVZju/7B/FA
ppx77Qmj1Oawkgp6vYt5kw8dR9ta5oYReL8YdFIrtriN8KygD8aL/THh5Vc65KXK
zd9WsttKj9AX/udwZ9SPT77uL/JehIQWlBY3lQhRPKISVr+PMfZQkg2ENf7xNdrF
vyFRBBQBDKjHVF7TCxOBIY7cmNPaHq1Bwgfjhw4ob7n+ncc79R9tTm/d8GcwVRCZ
ienZ9iU3g6lLi6FhF+/ku3PF/I8aa8w7k3U6cBqpeNkCs7GFYkkoH5ak8sMcN9VB
Lk/THRKicbn25keOKooZ9NofAKJBvQw8rf/7d182jCGZQf3T3Zw+jVTr9RIuJV6j
eXyIDsAedkXmcabmduwHu4QN+RG0OyqI6wVjATOaB1N3DEpFt5Srd0iFXcYhbTPd
pFQWjYrjSojzF4Un4NKR8nADAPITonPbGZBmQ4j8dk2D9nOiOajoJlR9BwCfZnUx
OIM4J/4kdaUqBcLXP3ydw9j1OLes1odoLO8iCFL2QtJ+sMrzb8DaCxQH7IdTcJOz
kb/8AFQfWijRNwZN4+CeTWo0rpd4m+jTO7ur9RyaEIRsUt25L98nseAc82LiNilF
yyhaC52OTsVbu/YZZZlOjBx+3UJflshdGbGZ2CMKB1ohxdRYbmD1/VIqO+lO+ICE
SgOsjRyfiLE5p2X7SpLKRqt7WvKDCzp4iBBDXqFMZ8i7gdaVaJ/124qS8YD2nwq/
iRYq0pMuIRj8Mzm+jetjgYcxwSH4xbdGd4SI4Kjb8VUX4zNYL26ckXItuk1KV/VH
u1Kli2B2UpnkrhmWlJ7S+DK0uO2V4PJYZaWHIFd0NVd12/xnt/9M+YriIvt9SoOZ
ysATRfAYv+UPcPhhmPVvQ7Geon4ftu09fvQZcpQztzHyGCE5JbknAHPIZWODW4kv
MnrUJsUHFW4Uz+MK3ZtKqfDGmU+kpNHCC1o3kRVt7Cz6eAcvUWrXbb+CQFmU0odc
9LzYBgwXmIgDg9FwSikdLfuDydKKtJCkddEefBCffjShwZCYIpugfoVsX841/6TD
NOpGfQMm+RDEkZWujDu7yznor1GfWGs2/9S1kQCz6mXfSuvY+Wi7Owtt1RaVvdGI
dkdSmJwF1/CZkqjGvtCZL1QQXhak1Qx1X+v9I7d0HsAyg9i04DM7Otsx0ftPDoFT
Uo26epEiqfyXHdDmw18etEi6cPRZztMXZ3yd5T1RUf7cFH69twYGbLjNMdNOGWuo
NM3UPtxmDtmIRSsr+RFbTwYiYYYp9END7fZkcz3TBtRk9MK0U62t4y1VxRnnHJ9N
XOAZxON5La6DMmVogYPNWffi/0GhO3pnpPENQXnlPLUiw90rSUeFcybIwOAb48WK
FzfsTIjpLKTRXxecrSdK+tFKXnbvalGbHTYMyWTJj1kKlQ1bkk+DIa1JtaKN4v0D
nnB/+HOYVHlu7EXPuqY1pZVMObubqDIhefb3EXOVInQDKSULzkjdLpFQ/vqrC4xS
H2HMWfOdR6VtXAqe6nhOpN+SFdxl6r1YxyNtp6P5ED8aRdE7ZWe+UPn8AjzxZjMS
TswuN02CweJ8aGvQgS3exAays2m3kQkaGqcaKJLjGztz+2VsKIwUxILS7trmpFcn
0w6hx/JRH+z5mwOfAZaY5k5ahPJSCZiNTFX6LjRqXFffOfl6MB2vpA5ifTHJvKYv
5HcrhLg2sklvsCxhAC76h7jtylVLx8Oap05WyX7lL8imgDnz4R4ibLUizzLkP5+g
39huny60o9A4XPLtEDcV5HIb5azEJfPg8FwBco8Supn9vYGam+QEvu7VRjYGLKVd
aBNjB1iio6p4mLh4b1PNm6/JunkKWvWLCD3GFX3mZuY55AZ2sx1gkXkxUABcvO8b
eAMTro53Ak4Ha2wvOFwsRIoJiLc0jYvQGt4xA0Vs+xdrKBVLrk/NM6eDSnKOXDXO
r2zraVTMZ/dcKGgz/VRa0Qn3AjI4B20vD4BfHCbNWUxVXFVIE/i/FMie+Netg0wg
PJGoYzxYlntArHyxbfC1WtcdtOrQYpmDUXHb5m4G4yE8oSIe2JTrRL36CkQ6g4id
gwjZEcqssH39blefWU5Ksd8B9GrtbY9LcFgufMu/7s1u3CRWSVlsfGgiuPP0CW8j
oYbQblWcPm1k1mM7R/5Kchf/sqkH09kpE/ATEXqThldZjK0BuRpTO+Bp+Lvxrvcs
dSt415bvATtIjiCcB+JIAXD0TN4HJgPMIBO7HpS5aP2Y7HdE0q3FyC4cTnUCz1kR
izEY2IZs5+UB+seUNSsw10f2qFBsdbAfJjHSFz2uLZqbYI7KzQ7eYv9TFYaQ61e6
O84cXwBVdSmHYFwFqMI7KLHDi1NftSzqT4GsbFoY5wt5aHULEJQYxv9S10msSI9O
HEthcm+QU3uUNwhsMU1cTcycvZD9t6ux4WO+fmLcvekMDsyBGELny2ldvcihQEeD
qfa76blYMCC9aJHju4GtQCgsc/18h3ovGhk1jSXBrCfbTBGXrnCgc4ZPrLlp/yPo
HCav6Vc3Ig792QEln5xOxVIGZnyFATZGKBtFvmodAZR41fUNA4G4FaFmtrLY72gT
CvE/RI8tfW4WJBL/Ch3GeBeUP8d/x83oaQ6JgbU0LL3+UkU9PVh5oy1knfjnSDUR
MgcBfvOPrP4/jMH6upwY/tlDQBpL3HnOcF/DrVbAxBIIAJGBFxS1bH/9XJZBcmg8
o+cqatukiwYHmJcFpVT32m4on6MxLBi23funfqcaddAkfSRUTMv0VPookI+p0z2a
CTZQmj6dukkBKdwNsnzO8QvRQplEPKzeHDKtvVcmaCRE+oWjCzQ19kSQ0++EhRd1
j14cOlVUQrHlt7N38m2WI8F68t7WnY2n0zQzsEDk8IurpEDaPH7+baUB+QcPQxwY
5BYcYdgFd7JhPwcVqTEu1xtMlPXwUjgeQrwRrLVmpuW+qf0DnHMfwJGSXDUAHlFQ
zeci6mSqpTwAv9l6gKAM9JrrmKM/BXztoixjy9AWkYZmcox9PEBlI54MlHkJV0dN
JF8+odj6fljYEzMt1gDI+C4a00nkVT+d1AJOYYa19QNjZu/K7CkUblfeUS40HhIm
pAEo39ujfAdsiT0I/LWzzdSEOfi4TpEWUy/QF9+FGdjecJ5FWfY736BpmPFOaL7c
jNSgjKNuSkWkIboL9ZCxFMoaco05TJWofSIgTJH9BcU3Fp5e+cQt5qcReY3Ai+Q0
fwaJbfVHz0+dhlfrgZaVoT+ACKSsitJrKaZaAYuvjrY8R0dLRTZ3xE9bIwXXEOrr
edM6+eoIR4LhPyga5QMYG4FWm8RZ1TjDYJM9rXp5jKozss/dArpE+hKImyOh+yHs
6MKo6O5cVsJ5ZhBUcTlxXpvWMpeRYmcA8l6GdCtBHTpSD6Ma8jAybOuxMaIzXS6v
nB6gT1DDqrqW3quEEEn5WV332FGyLF26ZRWMTQVsMRiR4b5ZFsKRFVVw53o6VlW0
LE6Jh2TRVS5KVBCzKBQkFgZ7j1MUZFbUmwtXh3fXH67UrgVYKg2YBR4AUv2Sixd7
Mrv0slf4wKIumzOY074LwnNYrd77Nm8vPAxfw+LegQTSaaXpJPCiqkCiEp6Fstw8
SBVWWecUBhEyJwuNdI7f+8I1ao2WtDXawPamkZrRSnA53hmEub6b2Xxzh9vHhbxM
AhfO0hzgh9DEI1FO4cq5x3e2b4SAwMUMvEk/9D7c3OBcF/zzLDcju3e/cpt39xyv
WvjxYx2iGq1Rr+55RZNfSXyJsh6C3VXGPjuPAng0JdsU1SRpKo8zFhAhHjkfl39K
qzV3vquLrITksZceP/lGIa8s5EBBFvR4n3ukeTYFGnOCv5kxE3MqVAqFOImwLxve
LYCPIzpvtsrkhvO8KVPicaL4yFEuIl/yeHvaaOaJqImJ3eZL3oLQUkMuGUeq9esh
ZG+6OpkbgQ6AC9ZdlnxJXVdcNfPD0wmFX8MJ20rWsPHqYogDG7EdQMj3p9UeJ89K
7nZJqZZ7urU6RTE+oAN8N/49fi+GhG4ayItqVuMqliTcnipnTqlADhRiOAWvL3aN
/fXoG889Ln4ntnsP2jLYKKgsfof64JGkeYWUUl7qnKXnGylPG7UFAj1DpJuE9oym
ZAwpHE3Q5xTI/teyx/zUpogBeHHgjKdk+sFv/Bw2/rh19RAJb1ZLFb4b3okmSO24
yQdNIhCGQRKjIxC8H9u0v6UsaeAXm3dkID1JPwxWejSQ8jGjw2klnKFXD9f/e9Xn
tiHuryjm6CDRAlJtm5OUc1VhfMwQsm86+8ThnYrhGYSvu8URZepRjV6Egn39z1jY
hwzTzOEZ0v+UdwiquhYZgNAgc2OFdGKQ+6mohNRXd7vZZ9wn0Qb9hMIcyQwxBEkf
jO0ibEobGbaz1HX7m4vAmk2nJofGzQZsMe7/mMhc5kVnSaMs287vghePgRzEda7B
yrnLzcbaK2TEnQ7o1mIirtnmVECpKrM50OMXi5JQrOV0RpVCpd5UnAqqJ8UIqzJ4
JimITgGQ8WjO2+48EGR700gnzeOKKNa+shLrincCCQ/3NpPSArxuZvw64ppIau9H
9S+McRNbSbxQop+PXhkt0QewrZj7dcT05VcLegmw0Ob+NtY2pDT71BhutqE9t3Ax
20+CxBwFdisGOhhqADkfJropqrlvwJoD89mGAXtbT7/qe0KhXSVWr5qtBd5Vyupm
ko2SK7Xk2bv92k/tlJKq7oBnNu2/LqE5ujm05+IaApwPoQIOQik6/4SnRVkjywrM
p+CLbBhXhdBqT0vYrOlDmswcMWpfLsAjE4KJF0Wq85fYsSXWOsfsNU9W3QklLJSr
Kzbk+Qw0i4mNf3gGwI9YgQ==

`pragma protect end_protected
