-- timer_14bit.vhd ------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- 14 bit timer
-- notification on 20, 1000 and 15000

-----------------------------------------------------------------------------

entity timer_14bit is
	port
	(
		clk				  : in 	std_logic;
		enable		  : in 	std_logic;
		clear_n		  : in 	std_logic;
		tim_3			  : out std_logic;
		tim_7			  : out std_logic;
		tim_20		  : out std_logic;
    tim_1000    : out std_logic;
    tim_15000		: out std_logic
	);
end timer_14bit;

-----------------------------------------------------------------------------

architecture rtl of timer_14bit is

  -- counter ----------------------------------------------------------------
  component counter_Nbit is
  	generic
  	(
  		N					: integer := 4
  	);
  	port
  	(
  		clk				: in 		std_logic;
  		enable		: in 		std_logic;
  		clear_n		: in 		std_logic;
  		rst_n			: in		std_logic;
  		cnt_out		: out 	std_logic_vector(N-1 downto 0)
  	);
  end component;

  -- internal signals ------------------------------------------------------
  signal cnt_out: std_logic_vector(13 downto 0);

  begin

    cnt: counter_Nbit generic map(14) port map(clk, enable, clear_n, '1', cnt_out);

		tim_3 		<= 	(cnt_out(0))			and (cnt_out(1)) 			and (not cnt_out(2)) 	and (not cnt_out(3)) 	and
              		(not cnt_out(4))	and (not cnt_out(5)) 	and (not cnt_out(6)) 	and (not cnt_out(7)) 	and
              		(not cnt_out(8)) 	and (not cnt_out(9)) 	and (not cnt_out(10)) and (not cnt_out(11)) and
              		(not cnt_out(12)) and (not cnt_out(13));

		tim_7 		<= 	(cnt_out(0))			and (cnt_out(1)) 			and (cnt_out(2)) 			and (not cnt_out(3)) 	and
									(not cnt_out(4)) 	and (not cnt_out(5)) 	and (not cnt_out(6)) 	and (not cnt_out(7)) 	and
									(not cnt_out(8)) 	and (not cnt_out(9)) 	and (not cnt_out(10)) and (not cnt_out(11)) and
									(not cnt_out(12)) and (not cnt_out(13));

    tim_20 		<= 	(not cnt_out(0))	and (not cnt_out(1)) 	and (cnt_out(2)) 			and (not cnt_out(3)) 	and
              		(cnt_out(4)) 			and (not cnt_out(5)) 	and (not cnt_out(6)) 	and (not cnt_out(7)) 	and
              		(not cnt_out(8)) 	and (not cnt_out(9)) 	and (not cnt_out(10)) and (not cnt_out(11)) and
              		(not cnt_out(12)) and (not cnt_out(13));

    tim_1000 	<= 	(not cnt_out(0)) 	and (not cnt_out(1)) 	and (not cnt_out(2)) 	and (cnt_out(3)) 			and
                	(not cnt_out(4)) 	and (cnt_out(5)) 			and (cnt_out(6)) 			and (cnt_out(7)) 			and
                	(cnt_out(8)) 			and (cnt_out(9)) 			and (not cnt_out(10)) and (not cnt_out(11)) and
                	(not cnt_out(12)) and (not cnt_out(13));

    tim_15000 <= 	(not cnt_out(0)) 	and (not cnt_out(1)) 	and (not cnt_out(2)) 	and (cnt_out(3)) 			and
                	(cnt_out(4)) 			and (not cnt_out(5)) 	and (not cnt_out(6)) 	and (cnt_out(7)) 			and
                	(not cnt_out(8)) 	and (cnt_out(9)) 			and (not cnt_out(10)) and (cnt_out(11)) 		and
                	(cnt_out(12)) 		and (cnt_out(13));

end rtl;

-----------------------------------------------------------------------------
