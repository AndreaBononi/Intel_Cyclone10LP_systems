-- blockram_system_v2_tb.vhd

-- Generated using ACDS version 22.1 917

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity blockram_system_v2_tb is
end entity blockram_system_v2_tb;

architecture rtl of blockram_system_v2_tb is
	component blockram_system_v2 is
		port (
			clk_clk         : in  std_logic                    := 'X';             -- clk
			leds_export     : out std_logic_vector(3 downto 0);                    -- export
			reset_reset_n   : in  std_logic                    := 'X';             -- reset_n
			switches_export : in  std_logic_vector(3 downto 0) := (others => 'X')  -- export
		);
	end component blockram_system_v2;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal blockram_system_v2_inst_clk_bfm_clk_clk       : std_logic; -- blockram_system_v2_inst_clk_bfm:clk -> [blockram_system_v2_inst:clk_clk, blockram_system_v2_inst_reset_bfm:clk]
	signal blockram_system_v2_inst_reset_bfm_reset_reset : std_logic; -- blockram_system_v2_inst_reset_bfm:reset -> blockram_system_v2_inst:reset_reset_n

begin

	blockram_system_v2_inst : component blockram_system_v2
		port map (
			clk_clk         => blockram_system_v2_inst_clk_bfm_clk_clk,       --      clk.clk
			leds_export     => open,                                          --     leds.export
			reset_reset_n   => blockram_system_v2_inst_reset_bfm_reset_reset, --    reset.reset_n
			switches_export => open                                           -- switches.export
		);

	blockram_system_v2_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => blockram_system_v2_inst_clk_bfm_clk_clk  -- clk.clk
		);

	blockram_system_v2_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => blockram_system_v2_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => blockram_system_v2_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of blockram_system_v2_tb
