`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h9vZLtcFFpGWYHDmAmRL92o+PnoDHYHFy6MBy4R4XE8UVwNYlGA0OyhiCUaP+gNs
SuuTf2ZJXnn/k6mNIs0gg/RRNKxL7qFWhAsSyH8neK+pSx57XvZ+2qs/Ause+a2p
BSyWWHi/H5OwofRLtYr7dOUMkjYo3DoDxdJqYNAxvUI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12336)
pV9IIZyExfkZyJ1HcfRETga+zsqiT8ipticPJaX5DU+Fe+p/ud4mU7aZ56TzWk/q
hhJbRxWZJNrjOinuZh601kyouJVvW0napA4fF3BYz7XcrvTFyYydBgRNMa0GO3lc
XD9xgOsGd5FEAPSz5lsz38FObnLO3Xb1o4WPGFuTLE4Y9q/jOgygsC3UcgeT46Q/
3eQXJB1JkzmxGOYwY3BeLmKrthlQnL2GwmrpyHTjrlthRWAc/s5xQhGVGhSSLTNP
AvrPIvyVv9nMZnfBmYXG0JyIWt99B76dU7Uf5hVAN7s84Z/9+3tUcz4/AUMKtLD2
voGk977+VMO8znPxnNAm8muyEf8POKHulfBSQEvjJS2rWXyvB7tllz+Aldz6YUbm
wQce2N47JKgGhn3MOrqcewzXQj7g8KHFxBbqEyTKZiEJPMMwfHnp815kDinCOKsT
RumURpnboNlO5joh1WdE+LQAz6/xm9rQ9+kf0IWVznFQN0LxIetE1BqBstOh8CTW
/Aboww3+0MPVHu0jEvbdwjrA2FQbjuf08/0EaAqy691OrZ6rv1JmYJPu9vvVhQ/V
96Keg1NfUT3GYgOzzHPHPRbERYi4k8vlIvqnbbb5/ySFK95FbFIwdB0KCRUHgkHz
nYusAUI/pjb3Cfro42kpbsnMs4yI+Yyn0fMNOwADEy5WI7CeW+AMahu1NGjTvemh
L8RBtfYUsp2CF2Cg1WG2fgIsjf2kEVyJ5xoslrHgBebyOxZ88IUlN0JyZVxpkAT+
kyrKYQN6sLNDi2f/KWkfHbK9wXgwSrkqWdD0imaS1l+3rMt3ws2hhiicoYU1Aif0
giYu5AOP0gTmwFrxxfSiJhPbgAPPgH3LLkNXYhdwdqO4pP+VNKcUB5klSJKTqYGC
kojl1w329A/DfPL2MO2HTYSbNdoTwrtKVK8atS5v1QdWLOq8t9OTQB3qW7lXWyI3
C9QwMVd8aVlwCT1R6cDkDygKWF17i8L+OCO/KQXv/qr89AI3uRC20tikDxUtzRlF
tT6CaQOWdq33h5IM0CYsZyEW05yBi/k2tQkZqhAu7RKNQT1FNs0fdSvjFHykHVhG
zycc/nQ00YJ9DUi1ETVbCdByDTmH+Mo0+0zlkdxOkJncMQptgqtrm7ZFyL2IuLpx
C0HCNDykHHMb0pSnGyJYzEStVjkJKHQ1NBKpf3A1+S56bZz3VzXMaWELynWYsInX
JH8SWDnxeGQrGH7itP5wADCI/sRy0hywTx0NlKZeWx2fSwqEynkeSiCB6iXA4CSN
/hyUK2iLZH/aeG1a3+1jHubiEIGOmyXnNJafofjYJQNV9HlsVaEFhc0KUlFoquRF
YfA6Ot4BAY9PviEsiiEZx7hWsWS21GAnBCW7kJooQf86K2VA9amr45X2DVgqSSid
qoQsug2ON8OYGHGuRLPiYV3zAhUI5Z6jo3juWhT4gOkvIm+moc7iyPl0ght6vtk2
q6CLQy79pUQ38SSKhq5PdkRg5LD8HAgwsPYN/1j94zuoC1Cv2QMgMrXUMR5jQwja
k1CmGxxA9VAhLmtnvgseiC6DKsP7tcD0UWgU2E7S+1/YqNogh0r85SBIPnG61g9f
jWVLI+SSLu3PP9QkyKq53ZRhfdepfDdXsQqk+kGFUIZjAUJC0gQTWh8FBbG2oD1T
y3YeFl+UENGJ9d8ifiNE2bA3oT0EVq+VKRCc+rCx+/3sp4s0Jksb7/fAOURfpcKL
AW1IwXBz3xmO4If/7zzkusPrTLT0iTRz9UB+6B3p8iayKyHoGt2C45G7xvRX6Xoz
I+NgMlDTTaiM9sr87dEenML70Zkr5qr/DJ38IucIHdfaji/AsaC86ny3mgVnRLaf
COC1kQ3OKNvQF0ebHC6Eo35HA4RlSpLK3B3ubiLMrfw3iwf1PBIndGmGOIj+0Xyn
NWvWijZ3yw4UTcGu/2jbd29IZQAINqz/cU9OP0a6J1QC5i8NqZ4ObI2J78mPqcuZ
XzV2ZLo3PQeqGT0oZEIC6RNCUGA975KOiN+1N/nDTYUiJiLyg2DYakqE8ogW0cK9
uKKJZGNZdok+yz2HP00a2ak85cAIhPIc9RqfgpMUf0kJN0SuI7FmHq8NNk/FPkmF
Tihv98uXUNpuVj/4R+VNn61sBAjw6CUSwAY6NJ3I8U4VegeToDaZEgH2B1eY750H
K3cYQmlNxnUsG7nE8O5rX5i3cGnhdKMCgFmrEWgtUq0drup+2Q3UyH7cd17TcycY
pyiGyPZ5nUZakdyImdlYcmyIwQxDusK/YkOL+PABuaus+n/u93Ri7+GBi+K3Gg7Z
f+fVb0wTrKDYV65l+78Moal1BNUTOqdKfbuCk0g2phZC/oT02VCdpFYbvyNDxoHR
J2z2uookByz8IQRKYrcCb/f/AhzSHRIujhG0+bBbtIQc6+CvMutyhEpM1z5v0J1g
2mliKN8YMh+wV6DNJhxiwxfBMtkntEyoNhnd//zPWCaT8qLcj0XW1fXJJjznnn9P
GkRWEJAry0bVJgv7G/HI2mr5FqRWAnFWsaXYdbFuGaHCVxivxmSggL5Z6bHX7IpE
NmxUw331ZLDYBppdnqvKL8SKEcDzHMbf3DFH6WG4Spq33r4tKnLqRtB3eTKMtJdW
3byCONneUIYLGDW+kk90N115DiEmIV7hAgZvrYabYOjjZMGhLvuOIxM+lnYgdBej
KZKTLxxOiLfj4dskQDkRu/HRhss/X4uFLrYc3XYfzYOnEm2hRHCaOD7E0JB85XgW
3DWqa56VISj7xlY4dPyjrOBdZS6tQSCOcFF/bE0tPbUDn+yd19B8rOZjJRQbMARp
Cn+zppQFc9nkv8VE2ZxkzPGPOI+W9KA3p2wIBYZ2NFzBMh8f7yB1x9qGww6keAIP
93yHldKpZ5hTPoZIlHAAcFiFxdA3wyAnu4in15MK87UMo1BSRBaMdmAisqxgWAXG
FZUjQtCEsZkyzi2f0xTgZzFx8vSQNV5kviBBb2+QPZGH96RXAv9tI7O8Ic//eq7H
ZUv+z//xi7JC5ZkuQrTtxvTg20MRtObkFGDErbg61Vf3eOxDZ+ygVXDsBmHhLxrr
NB0Im6Onwz1ds/HbW7WxjL+WNpRNMph9LwSmNsTd6qTFJNzgRFU3i/lGtAKmedMb
LcYThBKNjWXz7/kp18fZnFADbJoxO/dH/k0NL3cVy+YlZr6ccWaUH166MKfea76J
i0/Ku90uy0aSI2NcVyoZ4M7rHWGMAMNsqsVtHx1l5ZlxJOGhtZHnf/7Bo5cjFmy7
hE4mvYUFMzr1o9NPAuIifCNJ8O2wYhmNfwyXBiROSGneE6YCfiUKgKCUkf15yM1k
GZQ28H8KN5FB4dKrPLiG6X+JXrxLpnXEAgqBRoh6hvXSKvWNraOUv6pDagvN5rZQ
fbpIVLiTawK9UJvmBd++ojCDQ4uidnrL1uHSjg7CKlQhhf8Ha/biEgRZXGWUfM1q
YijjNFvKdiEM2pAhybof6fkI1QHsRHLN3UTcCeuVN4GhC4mKahpW3huc7WIq2PuQ
r5vTZ7mh7n+E7hacHJ7ZZKb+uDl8g9mjfQO9SYguXvEiC2/gFVkJfqYD8x8H9qSu
SjS2Df6o3FZdLXCJDG28nP7sRy2zPxlKkfhAncRXymvNEAPFad2jbmWAFMHvpDq9
KWmheSm0b+tyB+1G88rrDMStP7WX5BZZGxbsWka6GIeIO1xubtULx6PVn2Al6lNC
N0eNERdJ8COfQB4D2qTZwfIY3Hw4otFqSi1haFFk4KVEqOA7y59NmruSQTiGyfLb
cZ55AKkwxbXkZ1Regk6J9eepEpoSjI44M0j8aVGuhZ1qCQDOXvqcO6oqOv83ygqX
Rcs/Q2VNTHi7lRRHyoQ16vc50pqoU/4ABK52epCZg5LZfTmeP63u78GBQaB79esI
ob5pxvnlFuuiRW5nsvSSmfYudNDNUk/kwSc5ujo0t04STbIv0wYwNHhsAs02oH8m
pOqCieqqFmu82/LujGw68WQ3m1wbs9ErhSm7DPpELgK+aUtnBKAjf3qX406oy67E
tfHMOWdf+g/IQoaesBt5PJdxzQHOucdiO0cRcljTnObZNeaIGNa3U+sMjSvKddPO
tbJIw7m92Be6dwyjWrdSDdiH3J8VhX+QodJXeKb7XV7LjyFYQpS14ZFXQOjsOf2c
EBkSlK/i2ISZpt+GnbtxLfMwfCB5erih6PAhlTKFSen/9PwjVmwKdb6VMgbxU/nr
j9fUfhYTWEbWGysLE018O5WWnfJt/uvDPdH7Y/nJJVb4twbUw0en5prfuXrref2x
m2MwxkioXRqjGUlLFNw/rflnznfMTO/RHhiJ0Gp31/fJVytGjfVIDrN1HLIgeh1x
bh1NQoREVDf8WRq1XEI3KeV1Nk7NBPdE86+cHi+sWTe4PfiXad5S9SbpQuqFVK5j
DMmnf7qJPRP8rQJm+WbA6lbl5ibHGre/1tKg54Lv+fg94vcJmzR1G+k5DWjnkxQt
hqQekb8tMBSJx/pq+Tf4Uc+rm22lCk/NkIvGFdjTNT5ug7x4l0jsnAoDf5IaLmmz
cUnexfTOzo9CgqK9sqxB1WLihWMMPcRtt76N/SFB/wCw7HJmgE5NK1MdRCgoYIOO
auiDY499OfQv0KAl1930LjN8PaReDOMKvTWEAd51RtV9UCiEAOWi7tYqJMDK6Htd
ujAfNoDqLSfnpxx9wgv+1AIns5KWWcHEM9+0bMxesQa6YUVrvmGRQdaDwHXZZ/0C
9VUD2YunlOWU8+uTjepmeqma9ag+pmWTT3DO7xublbUwGRu6dyB+Cr4DOAfjhmcj
3rgWBtVtkVrUjWNEL23e54P9iP+nJQatpsA/VPl/XReSVTaW+lO06sbXrLNSx16E
RtrBg1f367G20K8yDN1+phUpclBplr4TKzEoFLeB/ELBhg0e02XtmHidkApaaPu2
8u7QOwEj4cCicXrhL8TK2WNJtVf1Vw3O+N9Oz8KIgrcebDT4cZLhStRJPOsHNFId
4nSjlf5MTn0yJC+dgwIOLyugcaGzSdlhIGxHNuw0kRqO3giOv2OMClm/BaCh6Cvw
rLZ41TCH76FMg1GUyANnrQmIbZoqYI7nUTtLqlLmR6nTPF7N9haNFaeCn/tTpDZI
Po5+22D6L7iC/GvmYUmHM/6LYFSxyZpAMCiFENouzxB4Dz5/SAqhEm6kDO12YBZV
EfZjVdaX6inAlNl2ogDMDyfuJUYIcKuYNx5Vtd45Tm3Qw3pPdUh2FxOboFFSXF06
pfQs/Q8xx98/hwWm3ZrKvJWJIikU91SWRtQgNXNBJ/D5sCCAIYsNqRO1iAvd6ePf
+hpDEwNpu5TgvLYOjJzsiBK80XcdU4v7k8H+FdxhF99cKUpZRBpz6SMhKPcgkYS3
PhKUocPIXFTJvUA9vwDUdVUes6bEE8AeHXSatgVx8nwFOYkTZGTwff0MQgXMxgNs
ztAexTYFP7TsbmKQ4jfRb30IklccNRso3NgMlJF8GOW0D/iXEX4wuuec5TerPntb
coFInFlDRs3HF2TalVFghKm+szPYYMx6OeNvJwAxiAJHtZHlgndybuGBIEi16qS2
RUn42LR82RNmFlSilGsSldM5Oop4TT2VUuV7KGQiyWSS8D25HyftWlmEjqRpi+0P
iR4sa7gyb8OwXrCChHOO9ULW9tFPf1GAtXEIrcGXUXEOiTzE/+EfgG+yDsO95IVm
4HXE0o0IbGDvdwGuIh0Z9MTHUW/oJgeZondGzvvY2aLPwYN/AAipagE6pgXvtiCM
O0yR31M8ylcycii+Q+nSW+//z0xc68aZwwB8EUsasrAq+1yQgLhPcy/nSs+5OQFd
YzNPoAN9wuBTdTaVD5r/ik8p77nsXqOIwCDlBzHKbUoyZtjh+akWMv6w4B+7NB3w
JUH1N14bPLf3/xRpj9oO7iRIrwhxyBell8rbXmQZguYTYVms6WBk4OGEc9eXi90r
/lUQQCcEMvw8HSUys22Ld3rVludPYXxM72MkP5TKZm7K4UrIBKtEmSInI5Zjre1s
ptpb4yx7YIahFMP/Dp7NehfDa+DaeBTOWbtp1rlYxiVE2j19VvdWFEihalsfAmC6
g6H1Mbs4NPvKUlqJooJqb99zn3RdBsZmq2ykR1So8tUSJAoq+Ul8V3B0f21OID+O
GTP5z4Rl+DK7mr4soCYn2/l3pcboD6I4JbLlQI+Wqw6OeAPGIviey71mhc+w9OjG
hGtdJhOiARdVr7qy4iRtV9glYo6EzGP/jUgB0t3txhnVZH58VcrCSR1q2cPUgBWo
MVi9tOMdcxgV56FdwPvtbF0PlNieyp71hIw8JhnR5Jjb4ughcz4surEv0hMr8evx
436xZO1HPxCrAyCVOBnWXSJW1JGONshfvBTwI6pIGImHD39mC6UZEpyZoUTi59PG
x5E6un8vAn+xOE/Kbk1Zpy2rEvGdOaTCK3cGK0Thhev33ybT8wmSHEJTgvrXv/OX
OE0zaT3T8tYNrxUAZNWXQJ0xd4cU+vyg7Bzm3n9xTQHCLJDv09cXi5/zTLr+vPQi
dlmsnIWZC8ZP/uQUCd5NO/l4ICwxKj59EVySWWcMsfmqDARvhlIZeB7cNybfo59X
s0cdOuZ4x8rGTYakZG8sj8PNeDGgGPLsgsFpBzPugyeHiu30O/EW0hwrUKACgNAW
7eZDlHzatnvnuwXasQMgI2L0srFTqVoUDRq6s7fWNuvaARQI2mddJzomwG6Gs+aB
/oHifQPSYROcQUc9yoHIswTB/ljcQnzPbj6qPYg7ot9OWwid0zlHg4BaDyNwBy7x
Rtg2iaVSwVNNSAchX+/PBxZVRpiJm5J9MrHYgiB0SBzt4jDh5BHbVHgM0+oP43ge
FSayyxDqiDveojNU5NkTwoqQApjnB7zT4SjTAfRZMpQuXyWKfkuWrs0I0ruSsLjk
ow9Zfd2EgkmS0T20806iow9GhSljkQh1mtfKrN3bfxokTjCHnH6391ngGGYPVwps
cZujBj4bg8So4xT6KbFeDk2lCRWAOJHtrOHrI2GIWdDhnm32RvIvXmEcvfzbYBTf
Hm5PfKrYgCWvCyP8SdAXR7Q15oC1+IhyykXyn3F7ZgR39/BEXetU49xxNsA6CUSv
QZgQKwleWuHOAlVB/AmKvwHP/FrRRR7FdQkmODMINTJqAQ9spr8Mm6lKWxGxCfO+
JRmZPifN7bbZB5RsB3FCx43e3fAgtTb4T8iXNpcAlpmw6TMBS0lt09lEQGWnCtkU
9GBs4qoaMykY5Efe11ZEE78vOR21NsjoDrUW4sT812eoIR9ugLEwMYFpxHQzASEu
qyZ9EAO66sw7yEOlqHk85Mr7VqpHuZ2oJc7w30xPtlYWhXBjUeG9+qBhRZRjeaWn
lnacrvCsk0kE0IG8W+wl8qAegOjnaue/FMCdLwAzkDB7lmT8BSeFxIOhLpOLuI8R
Oajic6A0WsWncCD/CK99fhOdpWRfMfXbZXN984RG1OUeU33abv7QeJPMLb1Lz9QI
72iKSns76yFN51jTbeh4SUNomYon6/Rwd4KYCX5WTnzjflBbfEXPy8HGJqCkTQ6J
oCZ2JlQ5hB1egk2F7CjQ+qXVuxXQaXTZ8nNYLMYJuKcKn1kRt9569W6fydn+AZ6L
W9Tut53NX18HSmTtElU7tmeniQRc0LxzZo3L+vpPIq9Ae7zJ32LQuV0U4qGgcmCa
3N1wCHqqXaIlQH+Sv3dllIM1GAYfZW552cv2zLzeMjy+44MQ6mEcedLzK8bbbI1v
YFJlQp/T6bO6Bame5/UVzgQbviJ+c7xStMHzbJ9RSATXWGfgkYXcIfBs400Uavna
T0qXa4GBtBzzoNqeDLKpeZGMOt53VzHK0SVqBPqQKNGtLr55rLabIVcVoKwpxSPF
LpzcgWz4sF1nab/YWB+mFpTlGcPbyKDVUEO7BL6hkeDH74Cy0acNwbwKeqfq5Jve
LOQlmh5neA3vJN5Nk1Lke8mVf+bU/iHnBkLuXwQl6TWy+1FCif/01Ay6rXEIae+O
B/BQ+2fCKw2q2utX3KtrDnD9W5iVgkDCzM2EQLTgzhlxeCA7ja9QRKYocGEAgIFn
WWeUEXsbco7ScJB9hd6xf9kc6dxmmt6tpL0cDM20FMtKIf/UA8UPKEJLSi/7s9xH
kuEhv/LBAOLkLITwAH7praU+fXT8g1WqXWo9sTR+m0FjxEDIsfcH6e69vCM2RApg
vtRNX66TDG3/N3LCO6yd+KuW9oQ6PM21xxDREiinjXjwNQG/5A6W5OAbxi97yjXS
Pn8syoyYRigxOyQwuWfOeLJ/kdz9HTfFk6mqnHtxzRPH7seehXOJDSSIAco6649S
a7+OivT3O8PLyREnGx9USZxOnFHyLkaHxLp7Zw8RSLB0onJ0WX1Nus6ZAFxcCYIV
R7Bt8eleOinfpxo4p0NjxVhmdy+lc+kcK5pJWBnXjZcSYxG9B0YM1VLJwRV1TLCh
MAImHp0D/grTb6uVv/kDgeX75xXDB7oLmkNOLT0sHm9ico58lEo7k6B1+KYBGx+w
ck4vQFAyux7r7ueFT7tsNt98IUb5wl/E1UU2jwY6A3Ry8GXte/LpoeW7ZGOXFYgw
dzd1TkPf7fjeDFej3X/n0oLhqzTI4cx65dHN+wmF0yb311jw+urKOEgWtsfIcyFk
ULNaiN8jGPoQvTvDcVp0ytlJfGcmOSVngnDsHBixJZdVTa5no0+tUZk42AE7RSF/
1nX1sG4iMFW6qZWguHd4b+PoOdXg0iOQqPS/gd5u9mQPo9SacSbl+MhDTfQxL6fW
RpwUdD4bcufiCliJt8iwSXS3crtyoDmSGcLUmobNa/5oO/tBoanHTXP4L0yapteM
wxgbu6sCut9oXsFPEunysMqLK15d/8plmToDRXjatmra8WD2ZnFs2IVZB0ZUESEE
FYz3qxFCjCA3bvpKxhLywIDXWzyJvzg/kzpxIA4LV3FGhAYqPHQd8PnQCFMdFCXs
/7Lb5VPSlJ4bQoMJLVTKh7dIzzBOuJ9GzSW4zorbBvQ1+mWCgeCniQ7sqLPHY+0W
QQdALbVlZsDv0LzGvYES8Ferwt+wZR552h3rVvMRU7/5flD04mYVAE+TF30C0jtQ
BF5+8vE75XgS0SCcxuMNBtIGzxveTC8OLrTp6qC3byDAciY8INeFZJgfdrriLS8x
/C9rwBvdDqEQdX/BJziqOT2FmZczh5wFSLYuAKZiiKBmE0s6NMgMYXohZBpB3ij5
tpZi5RmLTBrkJp6J8i+6Q6qDuiFYtYgch9qQOJk+zZRlnKJNiTLJMdelrbgOeF2S
KC/HzvTk1YQOdxbpiOz4ackrLY++ncoWm2y3IrIHpUexjF7XqgKG5mkVIgcS1yE3
R4G1pcPI24zxchK3m7+dU6nkneeLyZRCnDYJ78KH9ByXgkS/wMq61cjx22t8wBpN
MX2jlfVx1GJM9yAqgKmf6ZHcGQtsIn6230Uh7iLfy0BxS8mYTxQC4E/Lhfc5sA3x
xBvTClky1ZLa3MIFvF66mBs8ZSu3F9BVmoeHfRg5hHvybtGg7M0L5ZPfG5lTSYP7
Wjhv688Y8TglAjJL4iK2ZfkeBfe7NScqXPB5y+3zPrOLEzeiyLR+OADp16qPNcGn
DZ6XxiBUqX+6ZGIzaUn4Req8GkMKfMy/B1vp6aiEX65XJ4iUxlaxp5ynd5o7aUMR
buuC2eVf8LpYlDYJL/2ubKM99IIx36q2Qw4qXuolzZUIL0jb/9rU/rRTi381wdZb
KLWSd7XHCUwyD9HiYjxnxA3Wl6GBz+bbwk7OpsYjYANrfgLBk1WbeDCjV5ihacYR
xzx+GgFVCPaVp79miuza67mTUjnRJvpx8Cqvc30k3TEr1yWUwQPT5ZT/j2O76B04
iRmL5rFrGa/4JqSF7tAVzL8O2hNR2AjWHrI6xiMwlfrSFHFNB4eXR1OOcKZnXPk7
0NMR6FMsmkT59/lgbWzMg8VUJ/q8Sea5yuWzM/OrOcxiv6wEldlPHeTc5f1j5aHh
qeVyzMYANHkZ6+MldbsMx1VDMK5WUTbbS7lipRCCaDxNfnv+lXuWvxUZgjCQYSoH
NqgPTol7mQbnIfUIH7egLrTAxWwSiNI8K632fcyChPsWApmESv6fgClu80h8IqHn
diw4QYfQvPbHGqmAH3YPs1rK7Z2SYB+zNbH5EFWTYc40TBp0n8gveASRiflIS0Yg
HHwkJ4bvnJv6Mwpq8iAi/gDHMkMuKQBFmVwwvtx5GviAKGlUaM9ofzO5HabL5FAM
i55m6tUdGtQhhOuNz6ABhk635axpoyZwigTEJFsm3DqfrKQO5joySEoCnH6CeUz7
5RusxCUpG9CqgsXaN1QFrLeLXwo42SxM6wigtgDb01862cquArP7jahtsbfDlIvP
XqEWjg8FbY2tDGaF8wfTJ4t71BGWRNWzNHPGiTZWLKPvGjH26eomSy1GLiQZSkOm
Pi6pdJ3UhomYqS+4CG4/O3z/mdOdVcrHihOJyBYlyZuU/v+DrrBmAfZJaMiX0f4Q
SCtsyo+hFsi3iqJrdRXCrQjqoczNa2btOruyBhh3T7mtNiocMjNochs2QKIMLLUW
8Re80OQM1GRRjgXwapm2WbWBWgTh1J/zcJs5gNxSH9lIAOVabqXIX2q5M1tTWsP9
nFKMAFLYJz80Fv72tsSi5h83Um5xA7HTGwkJglJW55Ws9jv9GGRqlPpHMpCyY69F
jd8xT902rTIlRQCHmprAGsHUwWUCNFf9+NLl1NTfrNqcp81Zp+mOeCuZStsb8AO4
8LkfLyNsIqOtuD2g1HLCo2naDc7P0L+LX7SOt0jpORsbCKpBr4pZ4wULWhlMJasz
brwYSXZEtZ9iRe7ozZ7oxsi7hjpLMy/p8O+iNmWmsz17vOX0tr/qhKkqEDcyZSvk
tBRiVVwrDjeg/fDvgjWZYmQF7uE9tl68d/k+nt2f+IF/clyNHVTVRXCfUVZtdlvv
ewRyMwDC8Ufsx1iVrW+59APCm6Q5p6mkTFYewHF90pMsozqLzOQaK19d/rCIkGVM
yLgtu61nrTQWDsSmCDuE+reiBeGAeJJUdUASCYtDoesL+I6t1Ms7iotP6JTqwowK
4GW1mJIXspRPbwZFoQXIyXFE73OLT1j2mERj1PQjgxLnZAOR2SQPetU071ZhdIay
lScjqohFDn15Oy18T2kDv5Gl4IefKwHwHad9FNuWB3vw4fcCE8RmaWhKoO3wXkQx
WEvqAyIleteu9csehl7pJkecv9VXZLA14m/zugAr61jSkD2S3TMvzZSSvlVOMdyW
BUG+9IKfEWTEwa7Tp208OAqDRrarp9TlUeFYgXR9N9vwL8AVh5SPmzEJLdS9cFDU
qjgDR+laANezRvp461cMAq/SM19+raJCAZgOLE08xH9dBjhHqyeXI5T07TVBaO5P
XtWTlTlpuhmpu//GiKaF6TQUJqKAoWuWTpu4aYxz/NjIe2rhSbQ8TMhqqslf8Kh1
rNUYrstQt16/uQThJGhvE+x0bMmC7adH8B2axeoA7jvogKBhaJiIdoROWMtEHSpD
vHsj44EHGMiTO4ZJbJCMNwRl4lkoJh+udiTbdGS4FeX9VuP5yhFxNXJ9ooQDFYKa
EWcM79+GlUVTq8ju3reur/1wAaV2qeuncxKY7a//ioK76jtpbEQs/hhaQvQQ9W8N
PoORKh9Evrp2xs3EsFwRtLwVRKH+fdjCkRCDIHtezvffkeczi5i7gNv0UTQoFlZ5
KgYDJNvLV/byOvEj2zEmz2qayk74sjOHqx6m0mhnnITh3Lc90J5lpBYRXU9zXHKO
DQjuq4qOSw3dKVs3LfazmvRu48TNWDM7OwtBe1IY2GUgwrN/XYTSCH6wDlM6zKsX
oY9xXOf6H+zwoMDIJcwVIUZgex6ZwdhDQhvVlAr2VZhX4TI+6lv/LqUtvNtglYLU
EADt08A9yuWkw09NCc1ArlcCbBvlRnBYb+NKUQTIlmK6PRD/sRwKV2+4pIdQeoaq
cYD1G9GRuJlO1i6Q/2spLJrnz6cUvEYPmF3I4AyQvxWvgSJ1wMlMw8QG/iXTARWd
FfCz1KJ2ImXZxaStZIBBbfaxrVhZQbEJAFs8CRmlE8w837GXsJ8Lqmvat7B7ED4U
wdFt8yzFMYTQHmVHmGTyOgvtc9QUQtXcsLg7/QipfBmFs1h0c/DpLEmzumQgpIgk
IQUltpEkjqR1FkaQjVBfMj3ORnMbpWBjvr5aQCV48lCzgiSyV+yBYJgAhDZLVnbs
vlO5LYwOEvBZ3oUKb0s2vGrdryzo1LHfiMh5q9UvfFBhhiXWOsXVa0QAeFvQ14x+
b6wN1vUf3+b7UbZukvT8WwUTXacglBzHKmHVA8akRsU6LRZF/3ed8npeeuy/wk2r
4p56MRMQB/l5LIncSM7J/EluM20IR2msKuR4R428+uqZNgStsrd1E8gHhrkhi5VZ
dvbtjwSbUXktVVJ5de+YJCYgG0CGti5gWsjt/jJNQphaeb3AvKQkXN5CNvvMXX3Y
g3LPx9K9RH1KDwQ2OTl0hNgXlZNj9OvYtfT+VlhiMoQ6WlasP47dllNJazhhhXK5
6TChu3xJ+WB1kB4u+YWJZbNsIbnMypozT0d5AAoC3x5ew1fOOuO1A7XzDULEjA3Z
RGSdiMPxITMDcm7rn72QT4UktwtyxPstY/8xSge/K2rCHBNQRtPyPOrbMIKgp+gk
jgy9yXnQ73xK51ul3RyezV+KFoyWOuPaTf8IdKTtCU/cyVjyA+xTNebHEsNoN5KI
iIspGKHmRfw3H0Rh3Bsq7mgKzyYCuSb/hjawain8vbf0A89SW07/T0UPUGfpwlXx
Mj3JrcxqANNZiOHEvPYmLX64J1Pyvb5fQHJhpcfsN3NoaW4KOABjfIilO9ayLrge
UxVhAB2GQyz15B2feDLcIvcc7jmZ8iYxBwJiekpc4MZdaPNtcegoh/BtALonHh5+
U/PJSCs5lifFqtPSLqnnCV+5f8tf6BHZDSscq0i7B6ec5GNi4aSVL6VCzmgAm9YQ
1ngYE8k/vQmORRpTqk6ne4HGReYrEszdD+eFvasyD4tbkx7G/pzedOtPr94Rc4dT
ighz23rGIn7ZyLVCrpKE2CM7DO76c/e8s+9kkf8KU0A0lJUEMbh7cgRjm3V7X28e
yfUUCIez3HjEki/wxEx0RvFA/CwGmIQ7z/qtOXw29nW4qwF2Ld9V02oBtyHD41Fa
MQHx5VEWcNQlxHv+NI5hpz5u/ehc6I/frLEKNmDLjIw8lRtlV1XV664DcncAHVsb
cFC/YWL6rIDFMhp7f5eg+bTxbNEKbaBQZDJ+1iHHIN9R3fvPv35B5IsKqDbdm0u8
hBds3U+2FK50KZ26cGolj00SZM5eSe9W3M+gUfbii1XBHFof+uX8ViGPXVNBunP1
3g5XteFy0fYdvXY9S/gwVhJRjvQSQ86c52LllODoh9c+hN45rMMyJbRes6HLkgb5
c2IzbUu4VQDS0PnjXzZlZvfXe2bOdkiB8vxwpr7uwE/Sbxzpp4wiXO9b9z8aGaGI
6FsbhzpqW66jXt2Gz97//IypE5rVZRdvQMEvYUqNGZcAJWWVypAo7Dmj/2cc5h+Z
7c51laoWh2e8ThSNlk3IYkDiT3mi6jTuG0hmmduiVEVVSAof9AqF2deWn/8Spkgv
W0357cZh5zAZkMbA8EXud8Eb4boaFXaB+V2plW3Sal/33YO7IFHjJivlJo5F4ULY
7vSHDmsGX+rr3qxCF7M/ijTtCsiT+ZovjECMx0jndMwNWPOicHzMduxTNtuXVjKe
bAs9OVncRhC5SNlk+Nx0QUr+9pvjbv5HceOO0fHOnFQCl5PLHb0fIoOyN1asA6Lw
ENoqJDGad070w10qm/X5xjQEi0JP+43+s3SjR+0y24zFdU5yJGrX7HMXZ2xlJQOJ
1oiJnW7UK4HA1JbnQ/6AHuPxuBIAwvCu3Iij2W/Fb2s/FaBPlawTR0NZA71gabAc
Zpfpojnkqcg+vJMZfFytHqREZqOKBeaLLZ57I+/u7mo491ueDfLrNUHv1pIzQtfq
eBh9m8X+ehKPnkm15TvOVyzsvpuUAgvKSxQu1IV+41K6zUfRMNCAM7CaWBMxk6bb
d4c2xZgz6FbGTIPqqWE55zfBlWOjI/mZ141u57/qFpW0FJk/JxpGY0eiScUtyMJj
ukb2AWHNcyQHbYtutg7TUKUE35OVOfKrw35GUTTjJOIyP0RSQv0LMJAatxLvfDg5
eMt6NHqMNCl4dnEWZx9XHM/mX/+H691QJQ9b8mE3bKuHSrm8Yvyxj7M4j0uskPAP
WfbuETJXNDhtM0JTkbAupXm9A7Q6CwG+CP6dSjf0NRy/rY70HzmzV9/d8yD3vVMS
Egqt9Wh250+uG4qZqEuazmW3Cts2A97wxlzzzlXKJvh1uLAeubYJy8/50zoIOH5m
tGqLqyDYMCwrGL9qMAotd+YThK37Lbu7GvocwHeCc+GRNeONL6zaRkfnnSo4miCG
6TLYgBKs3Y8nRZ6OHCNEaAg4Gk3dDc04XRLRSoXOPnpYU3cWtATLZfxTIBjta49W
PyBem8UeMD0vBZkh2lVOsCIyBUZSdgq+ELk2gWaPX8Ua9asG4UKkWz+TiCzgcv0r
yn9awY6+mkTuzOpyfJ/ujlr6C/QlCkscJX4dPhVN3+mk6z7y/p/+1sSVRL/W13dK
FBOEnQwah/8yOkxu9G1HEHZ2ukYCpQhsY047qFNpEPMBAG8eOryoX5KkddWDvq+O
US80EVEXDdeRykYtvORt6MFah2mF3XUJa7m13CeszuK0/WrfQfPCNlksEYyz4wzt
e1v2L/F/qD+BCYoWctCJ4cr5H4tT6L/B3/yMVMFPH5OFG6hjwvUHKv4MEpDIfXvm
QZuuvtDz3ZjmvZlxrjRLN0bYRnX+D97S0EvzqJ8vtdYIGk4e6kYqbRAQ1M/L2op8
+qS2U8P+QCTQRVa2UTBkgmMKvQs+EYL1HkdOc9rKTxsLShFKLBCouVXv0dlBGUSC
j5avTLG/XEG2tk3oILmujGvdwg6v/WoMFLbT6ha2gCBw7cbzcTLFNcYXAZVf/ZGF
l663ECsZNQZlVHaucdFm7pti0jWyGXH5MskPX+d1iO6//2IZ2FRhviRDolE0vCqO
FIEijYlsdLVCXKmU1QZMKVwwYOufENm1bzKDuhbEG29I5/rLr/iOs3pzpsBR2u7b
W0cPWZQOQCWfwGImcM+IVB0ZekxW9deKNcqPLQUcSbAxTx55lpYqsIpWLcKH3L7t
24MBvGOR5pH2iPvjDus7x7aa7mZp08yPxemkc57Y/mnCroTd0owIi9EUfcKxWgVb
GoocB1cbL85oCH9cGCVX2QmHCBGSbQrKax4txLWPamstQa0+0pCXhIkbiK+FIe6q
BGvrLQGamwyo0ZWaliYueOez6Bzjo92Sl5Nh7R4jNpHGPyA3STnWK0RuzKzdnQiR
gyI+lIft+awK9CrNzMRwrZe3dP1pNBUALfTe7CUp2o/UfeeHALhS2NGGfHtmYjbs
48RdFhE2UtgR7/vf0FDdaT5o+gwWwMjk2lgiHtrYn8WuSQvP7vRtdvqGAy6zOzWQ
ZLzrm9YZHht0xOiMFW2sZGZM1wzTHFOgO28VZYO+cgCBZYeapEdGZbemEW6gyxUu
7qJxA62X/Wuh/QiLjCY/+UVhQlouiAWTQn6emg5ZeioHgdg40Avovq767gtUWJmV
z3NZWJVCxkCjFOB4rGB21+i+0dlYF7xrTNMP5GouuJfZOi36fs3r4Tkk8MsJx/qy
pH1GXB6sspXsqe485KgYDxIK6t0sg/yI4fSxKQTgzkl+iTXzbWJX/E2x4NshXc+b
cG4n8shpe9P0v5W6J7gQmrvnY7M8sJjEOKKXbEwaB+aourTU0Zy/UA1U87LtLlPP
7Nj458MaglKpgKBuwXYzuLr6NypGCqXZfJZ9NQB7kzhLu49x6a880KbND6W5T/kF
ZZ14umSTEZMmuHzhB1stFOIte7nuu5KRg4hapftMm9kSu5XyhD/exY6VjpNydN2S
jLFo3luiZhXNClE1QmnmjjCCeIT6K5txvOPUO61YXsJk5Ussz4KrcdZXe3qjkJFe
pTJSJjbwuzo5oS5Nv8r1yivb+S4gfr8UAqVPxK01eCJpkoLk6CC3NfoF7TigUv89
AaJaQORne03ttouDXZaygVkgJurEYjby9F+COQR+uFTbNfmkmPCh56e8tb/d/MIP
/4qI5S7brAk+R+ArirjijAZteEfDK8tK/DaYBveV/sAWm6n/9QvSjFZOs/h/RZa1
X4MsEPauL6rcwu7nnVdUNa3Yx6xdzovipN/yN+abtOSThiHdNL+NzdiDSWfDN30r
N8DCFeW/URytojBYUiBhcvO1q1BeXFF9FDTLUViJcAJgxxO9aKNvxkQsIgvQWuIP
16QAmI+5Yh5902G+9DDVTxyN6qE4cKi7HpLcRWG7vK+HmoBEb7BC/xZ5quHnVP9t
`pragma protect end_protected
