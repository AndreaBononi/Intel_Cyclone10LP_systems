-- blockram_system_v2.vhd

-- Generated using ACDS version 22.1 917

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity blockram_system_v2 is
	port (
		clk_clk         : in  std_logic                    := '0';             --      clk.clk
		leds_export     : out std_logic_vector(3 downto 0);                    --     leds.export
		reset_reset_n   : in  std_logic                    := '0';             --    reset.reset_n
		switches_export : in  std_logic_vector(3 downto 0) := (others => '0')  -- switches.export
	);
end entity blockram_system_v2;

architecture rtl of blockram_system_v2 is
	component custom_OCRAM is
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset_n                : in  std_logic                     := 'X';             -- reset_n
			avs_address            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avs_read               : in  std_logic                     := 'X';             -- read
			avs_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			avs_write              : in  std_logic                     := 'X';             -- write
			avs_writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_waitrequest        : out std_logic;                                        -- waitrequest
			avs_readdatavalid      : out std_logic;                                        -- readdatavalid
			avs_beginbursttransfer : in  std_logic                     := 'X';             -- beginbursttransfer
			avs_burstcount         : in  std_logic_vector(10 downto 0) := (others => 'X')  -- burstcount
		);
	end component custom_OCRAM;

	component blockram_system_v2_instruction_OCROM is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			debugaccess : in  std_logic                     := 'X';             -- debugaccess
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component blockram_system_v2_instruction_OCROM;

	component blockram_system_v2_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component blockram_system_v2_leds;

	component blockram_system_v2_nios2f is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(13 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(12 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component blockram_system_v2_nios2f;

	component blockram_system_v2_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component blockram_system_v2_switches;

	component blockram_system_v2_mm_interconnect_0 is
		port (
			clk_100MHz_clk_clk                         : in  std_logic                     := 'X';             -- clk
			nios2f_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			nios2f_data_master_address                 : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			nios2f_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2f_data_master_burstcount              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			nios2f_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2f_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2f_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2f_data_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			nios2f_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2f_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2f_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2f_instruction_master_address          : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			nios2f_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2f_instruction_master_burstcount       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			nios2f_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2f_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			nios2f_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			data_OCRAM_avalon_slave_address            : out std_logic_vector(7 downto 0);                     -- address
			data_OCRAM_avalon_slave_write              : out std_logic;                                        -- write
			data_OCRAM_avalon_slave_read               : out std_logic;                                        -- read
			data_OCRAM_avalon_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			data_OCRAM_avalon_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			data_OCRAM_avalon_slave_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			data_OCRAM_avalon_slave_burstcount         : out std_logic_vector(10 downto 0);                    -- burstcount
			data_OCRAM_avalon_slave_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			data_OCRAM_avalon_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			instruction_OCROM_s1_address               : out std_logic_vector(9 downto 0);                     -- address
			instruction_OCROM_s1_write                 : out std_logic;                                        -- write
			instruction_OCROM_s1_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			instruction_OCROM_s1_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			instruction_OCROM_s1_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			instruction_OCROM_s1_chipselect            : out std_logic;                                        -- chipselect
			instruction_OCROM_s1_clken                 : out std_logic;                                        -- clken
			instruction_OCROM_s1_debugaccess           : out std_logic;                                        -- debugaccess
			leds_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                              : out std_logic;                                        -- write
			leds_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                         : out std_logic;                                        -- chipselect
			nios2f_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			nios2f_debug_mem_slave_write               : out std_logic;                                        -- write
			nios2f_debug_mem_slave_read                : out std_logic;                                        -- read
			nios2f_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2f_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			nios2f_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2f_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			nios2f_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			switches_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component blockram_system_v2_mm_interconnect_0;

	component blockram_system_v2_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component blockram_system_v2_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2f_data_master_readdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2f_data_master_readdata -> nios2f:d_readdata
	signal nios2f_data_master_waitrequest                               : std_logic;                     -- mm_interconnect_0:nios2f_data_master_waitrequest -> nios2f:d_waitrequest
	signal nios2f_data_master_debugaccess                               : std_logic;                     -- nios2f:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2f_data_master_debugaccess
	signal nios2f_data_master_address                                   : std_logic_vector(13 downto 0); -- nios2f:d_address -> mm_interconnect_0:nios2f_data_master_address
	signal nios2f_data_master_byteenable                                : std_logic_vector(3 downto 0);  -- nios2f:d_byteenable -> mm_interconnect_0:nios2f_data_master_byteenable
	signal nios2f_data_master_read                                      : std_logic;                     -- nios2f:d_read -> mm_interconnect_0:nios2f_data_master_read
	signal nios2f_data_master_readdatavalid                             : std_logic;                     -- mm_interconnect_0:nios2f_data_master_readdatavalid -> nios2f:d_readdatavalid
	signal nios2f_data_master_write                                     : std_logic;                     -- nios2f:d_write -> mm_interconnect_0:nios2f_data_master_write
	signal nios2f_data_master_writedata                                 : std_logic_vector(31 downto 0); -- nios2f:d_writedata -> mm_interconnect_0:nios2f_data_master_writedata
	signal nios2f_data_master_burstcount                                : std_logic_vector(3 downto 0);  -- nios2f:d_burstcount -> mm_interconnect_0:nios2f_data_master_burstcount
	signal nios2f_instruction_master_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2f_instruction_master_readdata -> nios2f:i_readdata
	signal nios2f_instruction_master_waitrequest                        : std_logic;                     -- mm_interconnect_0:nios2f_instruction_master_waitrequest -> nios2f:i_waitrequest
	signal nios2f_instruction_master_address                            : std_logic_vector(12 downto 0); -- nios2f:i_address -> mm_interconnect_0:nios2f_instruction_master_address
	signal nios2f_instruction_master_read                               : std_logic;                     -- nios2f:i_read -> mm_interconnect_0:nios2f_instruction_master_read
	signal nios2f_instruction_master_readdatavalid                      : std_logic;                     -- mm_interconnect_0:nios2f_instruction_master_readdatavalid -> nios2f:i_readdatavalid
	signal nios2f_instruction_master_burstcount                         : std_logic_vector(3 downto 0);  -- nios2f:i_burstcount -> mm_interconnect_0:nios2f_instruction_master_burstcount
	signal mm_interconnect_0_data_ocram_avalon_slave_beginbursttransfer : std_logic;                     -- mm_interconnect_0:data_OCRAM_avalon_slave_beginbursttransfer -> data_OCRAM:avs_beginbursttransfer
	signal mm_interconnect_0_data_ocram_avalon_slave_readdata           : std_logic_vector(31 downto 0); -- data_OCRAM:avs_readdata -> mm_interconnect_0:data_OCRAM_avalon_slave_readdata
	signal mm_interconnect_0_data_ocram_avalon_slave_waitrequest        : std_logic;                     -- data_OCRAM:avs_waitrequest -> mm_interconnect_0:data_OCRAM_avalon_slave_waitrequest
	signal mm_interconnect_0_data_ocram_avalon_slave_address            : std_logic_vector(7 downto 0);  -- mm_interconnect_0:data_OCRAM_avalon_slave_address -> data_OCRAM:avs_address
	signal mm_interconnect_0_data_ocram_avalon_slave_read               : std_logic;                     -- mm_interconnect_0:data_OCRAM_avalon_slave_read -> data_OCRAM:avs_read
	signal mm_interconnect_0_data_ocram_avalon_slave_readdatavalid      : std_logic;                     -- data_OCRAM:avs_readdatavalid -> mm_interconnect_0:data_OCRAM_avalon_slave_readdatavalid
	signal mm_interconnect_0_data_ocram_avalon_slave_write              : std_logic;                     -- mm_interconnect_0:data_OCRAM_avalon_slave_write -> data_OCRAM:avs_write
	signal mm_interconnect_0_data_ocram_avalon_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:data_OCRAM_avalon_slave_writedata -> data_OCRAM:avs_writedata
	signal mm_interconnect_0_data_ocram_avalon_slave_burstcount         : std_logic_vector(10 downto 0); -- mm_interconnect_0:data_OCRAM_avalon_slave_burstcount -> data_OCRAM:avs_burstcount
	signal mm_interconnect_0_nios2f_debug_mem_slave_readdata            : std_logic_vector(31 downto 0); -- nios2f:debug_mem_slave_readdata -> mm_interconnect_0:nios2f_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2f_debug_mem_slave_waitrequest         : std_logic;                     -- nios2f:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2f_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2f_debug_mem_slave_debugaccess         : std_logic;                     -- mm_interconnect_0:nios2f_debug_mem_slave_debugaccess -> nios2f:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2f_debug_mem_slave_address             : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2f_debug_mem_slave_address -> nios2f:debug_mem_slave_address
	signal mm_interconnect_0_nios2f_debug_mem_slave_read                : std_logic;                     -- mm_interconnect_0:nios2f_debug_mem_slave_read -> nios2f:debug_mem_slave_read
	signal mm_interconnect_0_nios2f_debug_mem_slave_byteenable          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2f_debug_mem_slave_byteenable -> nios2f:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2f_debug_mem_slave_write               : std_logic;                     -- mm_interconnect_0:nios2f_debug_mem_slave_write -> nios2f:debug_mem_slave_write
	signal mm_interconnect_0_nios2f_debug_mem_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2f_debug_mem_slave_writedata -> nios2f:debug_mem_slave_writedata
	signal mm_interconnect_0_switches_s1_readdata                       : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_0:switches_s1_readdata
	signal mm_interconnect_0_switches_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switches_s1_address -> switches:address
	signal mm_interconnect_0_leds_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                           : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                              : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_instruction_ocrom_s1_chipselect            : std_logic;                     -- mm_interconnect_0:instruction_OCROM_s1_chipselect -> instruction_OCROM:chipselect
	signal mm_interconnect_0_instruction_ocrom_s1_readdata              : std_logic_vector(31 downto 0); -- instruction_OCROM:readdata -> mm_interconnect_0:instruction_OCROM_s1_readdata
	signal mm_interconnect_0_instruction_ocrom_s1_debugaccess           : std_logic;                     -- mm_interconnect_0:instruction_OCROM_s1_debugaccess -> instruction_OCROM:debugaccess
	signal mm_interconnect_0_instruction_ocrom_s1_address               : std_logic_vector(9 downto 0);  -- mm_interconnect_0:instruction_OCROM_s1_address -> instruction_OCROM:address
	signal mm_interconnect_0_instruction_ocrom_s1_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:instruction_OCROM_s1_byteenable -> instruction_OCROM:byteenable
	signal mm_interconnect_0_instruction_ocrom_s1_write                 : std_logic;                     -- mm_interconnect_0:instruction_OCROM_s1_write -> instruction_OCROM:write
	signal mm_interconnect_0_instruction_ocrom_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:instruction_OCROM_s1_writedata -> instruction_OCROM:writedata
	signal mm_interconnect_0_instruction_ocrom_s1_clken                 : std_logic;                     -- mm_interconnect_0:instruction_OCROM_s1_clken -> instruction_OCROM:clken
	signal nios2f_irq_irq                                               : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2f:irq
	signal rst_controller_reset_out_reset                               : std_logic;                     -- rst_controller:reset_out -> [instruction_OCROM:reset, irq_mapper:reset, mm_interconnect_0:nios2f_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                           : std_logic;                     -- rst_controller:reset_req -> [instruction_OCROM:reset_req, nios2f:reset_req, rst_translator:reset_req_in]
	signal nios2f_debug_reset_request_reset                             : std_logic;                     -- nios2f:debug_reset_request -> rst_controller:reset_in1
	signal reset_reset_n_ports_inv                                      : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_leds_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal rst_controller_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_reset_out_reset:inv -> [data_OCRAM:reset_n, leds:reset_n, nios2f:reset_n, switches:reset_n]

begin

	data_ocram : component custom_OCRAM
		port map (
			clk                    => clk_clk,                                                      --        clock.clk
			reset_n                => rst_controller_reset_out_reset_ports_inv,                     --        reset.reset_n
			avs_address            => mm_interconnect_0_data_ocram_avalon_slave_address,            -- avalon_slave.address
			avs_read               => mm_interconnect_0_data_ocram_avalon_slave_read,               --             .read
			avs_readdata           => mm_interconnect_0_data_ocram_avalon_slave_readdata,           --             .readdata
			avs_write              => mm_interconnect_0_data_ocram_avalon_slave_write,              --             .write
			avs_writedata          => mm_interconnect_0_data_ocram_avalon_slave_writedata,          --             .writedata
			avs_waitrequest        => mm_interconnect_0_data_ocram_avalon_slave_waitrequest,        --             .waitrequest
			avs_readdatavalid      => mm_interconnect_0_data_ocram_avalon_slave_readdatavalid,      --             .readdatavalid
			avs_beginbursttransfer => mm_interconnect_0_data_ocram_avalon_slave_beginbursttransfer, --             .beginbursttransfer
			avs_burstcount         => mm_interconnect_0_data_ocram_avalon_slave_burstcount          --             .burstcount
		);

	instruction_ocrom : component blockram_system_v2_instruction_OCROM
		port map (
			clk         => clk_clk,                                            --   clk1.clk
			address     => mm_interconnect_0_instruction_ocrom_s1_address,     --     s1.address
			debugaccess => mm_interconnect_0_instruction_ocrom_s1_debugaccess, --       .debugaccess
			clken       => mm_interconnect_0_instruction_ocrom_s1_clken,       --       .clken
			chipselect  => mm_interconnect_0_instruction_ocrom_s1_chipselect,  --       .chipselect
			write       => mm_interconnect_0_instruction_ocrom_s1_write,       --       .write
			readdata    => mm_interconnect_0_instruction_ocrom_s1_readdata,    --       .readdata
			writedata   => mm_interconnect_0_instruction_ocrom_s1_writedata,   --       .writedata
			byteenable  => mm_interconnect_0_instruction_ocrom_s1_byteenable,  --       .byteenable
			reset       => rst_controller_reset_out_reset,                     -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,                 --       .reset_req
			freeze      => '0'                                                 -- (terminated)
		);

	leds : component blockram_system_v2_leds
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_export                                -- external_connection.export
		);

	nios2f : component blockram_system_v2_nios2f
		port map (
			clk                                 => clk_clk,                                              --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                   --                          .reset_req
			d_address                           => nios2f_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2f_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2f_data_master_read,                              --                          .read
			d_readdata                          => nios2f_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2f_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2f_data_master_write,                             --                          .write
			d_writedata                         => nios2f_data_master_writedata,                         --                          .writedata
			d_burstcount                        => nios2f_data_master_burstcount,                        --                          .burstcount
			d_readdatavalid                     => nios2f_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2f_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2f_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2f_instruction_master_read,                       --                          .read
			i_readdata                          => nios2f_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2f_instruction_master_waitrequest,                --                          .waitrequest
			i_burstcount                        => nios2f_instruction_master_burstcount,                 --                          .burstcount
			i_readdatavalid                     => nios2f_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2f_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2f_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2f_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2f_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2f_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2f_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2f_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2f_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2f_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2f_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                  -- custom_instruction_master.readra
		);

	switches : component blockram_system_v2_switches
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switches_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_switches_s1_readdata,   --                    .readdata
			in_port  => switches_export                           -- external_connection.export
		);

	mm_interconnect_0 : component blockram_system_v2_mm_interconnect_0
		port map (
			clk_100MHz_clk_clk                         => clk_clk,                                                      --                     clk_100MHz_clk.clk
			nios2f_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                               -- nios2f_reset_reset_bridge_in_reset.reset
			nios2f_data_master_address                 => nios2f_data_master_address,                                   --                 nios2f_data_master.address
			nios2f_data_master_waitrequest             => nios2f_data_master_waitrequest,                               --                                   .waitrequest
			nios2f_data_master_burstcount              => nios2f_data_master_burstcount,                                --                                   .burstcount
			nios2f_data_master_byteenable              => nios2f_data_master_byteenable,                                --                                   .byteenable
			nios2f_data_master_read                    => nios2f_data_master_read,                                      --                                   .read
			nios2f_data_master_readdata                => nios2f_data_master_readdata,                                  --                                   .readdata
			nios2f_data_master_readdatavalid           => nios2f_data_master_readdatavalid,                             --                                   .readdatavalid
			nios2f_data_master_write                   => nios2f_data_master_write,                                     --                                   .write
			nios2f_data_master_writedata               => nios2f_data_master_writedata,                                 --                                   .writedata
			nios2f_data_master_debugaccess             => nios2f_data_master_debugaccess,                               --                                   .debugaccess
			nios2f_instruction_master_address          => nios2f_instruction_master_address,                            --          nios2f_instruction_master.address
			nios2f_instruction_master_waitrequest      => nios2f_instruction_master_waitrequest,                        --                                   .waitrequest
			nios2f_instruction_master_burstcount       => nios2f_instruction_master_burstcount,                         --                                   .burstcount
			nios2f_instruction_master_read             => nios2f_instruction_master_read,                               --                                   .read
			nios2f_instruction_master_readdata         => nios2f_instruction_master_readdata,                           --                                   .readdata
			nios2f_instruction_master_readdatavalid    => nios2f_instruction_master_readdatavalid,                      --                                   .readdatavalid
			data_OCRAM_avalon_slave_address            => mm_interconnect_0_data_ocram_avalon_slave_address,            --            data_OCRAM_avalon_slave.address
			data_OCRAM_avalon_slave_write              => mm_interconnect_0_data_ocram_avalon_slave_write,              --                                   .write
			data_OCRAM_avalon_slave_read               => mm_interconnect_0_data_ocram_avalon_slave_read,               --                                   .read
			data_OCRAM_avalon_slave_readdata           => mm_interconnect_0_data_ocram_avalon_slave_readdata,           --                                   .readdata
			data_OCRAM_avalon_slave_writedata          => mm_interconnect_0_data_ocram_avalon_slave_writedata,          --                                   .writedata
			data_OCRAM_avalon_slave_beginbursttransfer => mm_interconnect_0_data_ocram_avalon_slave_beginbursttransfer, --                                   .beginbursttransfer
			data_OCRAM_avalon_slave_burstcount         => mm_interconnect_0_data_ocram_avalon_slave_burstcount,         --                                   .burstcount
			data_OCRAM_avalon_slave_readdatavalid      => mm_interconnect_0_data_ocram_avalon_slave_readdatavalid,      --                                   .readdatavalid
			data_OCRAM_avalon_slave_waitrequest        => mm_interconnect_0_data_ocram_avalon_slave_waitrequest,        --                                   .waitrequest
			instruction_OCROM_s1_address               => mm_interconnect_0_instruction_ocrom_s1_address,               --               instruction_OCROM_s1.address
			instruction_OCROM_s1_write                 => mm_interconnect_0_instruction_ocrom_s1_write,                 --                                   .write
			instruction_OCROM_s1_readdata              => mm_interconnect_0_instruction_ocrom_s1_readdata,              --                                   .readdata
			instruction_OCROM_s1_writedata             => mm_interconnect_0_instruction_ocrom_s1_writedata,             --                                   .writedata
			instruction_OCROM_s1_byteenable            => mm_interconnect_0_instruction_ocrom_s1_byteenable,            --                                   .byteenable
			instruction_OCROM_s1_chipselect            => mm_interconnect_0_instruction_ocrom_s1_chipselect,            --                                   .chipselect
			instruction_OCROM_s1_clken                 => mm_interconnect_0_instruction_ocrom_s1_clken,                 --                                   .clken
			instruction_OCROM_s1_debugaccess           => mm_interconnect_0_instruction_ocrom_s1_debugaccess,           --                                   .debugaccess
			leds_s1_address                            => mm_interconnect_0_leds_s1_address,                            --                            leds_s1.address
			leds_s1_write                              => mm_interconnect_0_leds_s1_write,                              --                                   .write
			leds_s1_readdata                           => mm_interconnect_0_leds_s1_readdata,                           --                                   .readdata
			leds_s1_writedata                          => mm_interconnect_0_leds_s1_writedata,                          --                                   .writedata
			leds_s1_chipselect                         => mm_interconnect_0_leds_s1_chipselect,                         --                                   .chipselect
			nios2f_debug_mem_slave_address             => mm_interconnect_0_nios2f_debug_mem_slave_address,             --             nios2f_debug_mem_slave.address
			nios2f_debug_mem_slave_write               => mm_interconnect_0_nios2f_debug_mem_slave_write,               --                                   .write
			nios2f_debug_mem_slave_read                => mm_interconnect_0_nios2f_debug_mem_slave_read,                --                                   .read
			nios2f_debug_mem_slave_readdata            => mm_interconnect_0_nios2f_debug_mem_slave_readdata,            --                                   .readdata
			nios2f_debug_mem_slave_writedata           => mm_interconnect_0_nios2f_debug_mem_slave_writedata,           --                                   .writedata
			nios2f_debug_mem_slave_byteenable          => mm_interconnect_0_nios2f_debug_mem_slave_byteenable,          --                                   .byteenable
			nios2f_debug_mem_slave_waitrequest         => mm_interconnect_0_nios2f_debug_mem_slave_waitrequest,         --                                   .waitrequest
			nios2f_debug_mem_slave_debugaccess         => mm_interconnect_0_nios2f_debug_mem_slave_debugaccess,         --                                   .debugaccess
			switches_s1_address                        => mm_interconnect_0_switches_s1_address,                        --                        switches_s1.address
			switches_s1_readdata                       => mm_interconnect_0_switches_s1_readdata                        --                                   .readdata
		);

	irq_mapper : component blockram_system_v2_irq_mapper
		port map (
			clk        => clk_clk,                        --       clk.clk
			reset      => rst_controller_reset_out_reset, -- clk_reset.reset
			sender_irq => nios2f_irq_irq                  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios2f_debug_reset_request_reset,   -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of blockram_system_v2
