-- basic_system_tb.vhd

-- Generated using ACDS version 22.1 917

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity basic_system_tb is
end entity basic_system_tb;

architecture rtl of basic_system_tb is
	component basic_system is
		port (
			clk_clk           : in  std_logic                    := 'X';             -- clk
			leds_export       : out std_logic_vector(3 downto 0);                    -- export
			reset_reset_n     : in  std_logic                    := 'X';             -- reset_n
			rst_switch_export : in  std_logic                    := 'X';             -- export
			switches_export   : in  std_logic_vector(3 downto 0) := (others => 'X')  -- export
		);
	end component basic_system;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal basic_system_inst_clk_bfm_clk_clk       : std_logic; -- basic_system_inst_clk_bfm:clk -> [basic_system_inst:clk_clk, basic_system_inst_reset_bfm:clk]
	signal basic_system_inst_reset_bfm_reset_reset : std_logic; -- basic_system_inst_reset_bfm:reset -> basic_system_inst:reset_reset_n

begin

	basic_system_inst : component basic_system
		port map (
			clk_clk           => basic_system_inst_clk_bfm_clk_clk,       --        clk.clk
			leds_export       => open,                                    --       leds.export
			reset_reset_n     => basic_system_inst_reset_bfm_reset_reset, --      reset.reset_n
			rst_switch_export => open,                                    -- rst_switch.export
			switches_export   => open                                     --   switches.export
		);

	basic_system_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 100000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => basic_system_inst_clk_bfm_clk_clk  -- clk.clk
		);

	basic_system_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => basic_system_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => basic_system_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of basic_system_tb
